`timescale 10ps / 1fs

module sys_test();

parameter EC_BASE_FIELD_WIDTH = 377;
parameter EC_SCALAR_FIELD_WIDTH = 253; 
parameter ADDR_WIDTH = 8;
parameter MEM_SIZE = 256;
parameter CLK_PERIOD = 100;

    reg ap_clk, ap_rst, ap_start;
    wire ap_done, ap_idle, ap_ready;

    wire [EC_BASE_FIELD_WIDTH - 1:0] P_arr_x_q0, P_arr_x_q1;
    wire [EC_BASE_FIELD_WIDTH - 1:0] P_arr_x_d0, P_arr_x_d1;
    wire P_arr_x_we0, P_arr_x_we1;
    wire [ADDR_WIDTH-1:0] P_arr_x_address0, P_arr_x_address1;
    
    wire [EC_BASE_FIELD_WIDTH - 1:0] P_arr_y_q0, P_arr_y_q1;
    wire [EC_BASE_FIELD_WIDTH - 1:0] P_arr_y_d0, P_arr_y_d1;
    wire P_arr_y_we0, P_arr_y_we1;
    wire [ADDR_WIDTH-1:0] P_arr_y_address0, P_arr_y_address1;
    
    wire [EC_BASE_FIELD_WIDTH - 1:0] P_arr_z_q0, P_arr_z_q1;
    wire [EC_BASE_FIELD_WIDTH - 1:0] P_arr_z_d0, P_arr_z_d1;
    wire P_arr_z_we0, P_arr_z_we1;
    wire [ADDR_WIDTH-1:0] P_arr_z_address0, P_arr_z_address1;
    
    wire [EC_SCALAR_FIELD_WIDTH - 1:0] K_arr_q0, K_arr_q1;
    wire [EC_SCALAR_FIELD_WIDTH - 1:0] K_arr_d0, K_arr_d1;
    wire K_arr_we0, K_arr_we1;
    wire [ADDR_WIDTH-1:0] K_arr_address0, K_arr_address1;

    wire  [14:0] total_num_padd_ops;

    reg [14:0] cnt_bucket_chunks_0 [0:63];
    reg [14:0] cnt_bucket_chunks_1 [0:63];
    reg [14:0] cnt_bucket_chunks_2 [0:63];
    reg [14:0] cnt_bucket_chunks_3 [0:63];
    reg [14:0] cnt_bucket_chunks_4 [0:63];
    reg [14:0] cnt_bucket_chunks_5 [0:63];
    reg [14:0] cnt_bucket_chunks_6 [0:63];
    reg [14:0] cnt_bucket_chunks_7 [0:63];
    reg [14:0] cnt_bucket_chunks_8 [0:63];
    reg [14:0] cnt_bucket_chunks_9 [0:63];
    reg [14:0] cnt_bucket_chunks_10 [0:63];
    reg [14:0] cnt_bucket_chunks_11 [0:63];
    reg [14:0] cnt_bucket_chunks_12 [0:63];
    reg [14:0] cnt_bucket_chunks_13 [0:63];
    reg [14:0] cnt_bucket_chunks_14 [0:63];
    reg [14:0] cnt_bucket_chunks_15 [0:63];
    reg [14:0] cnt_bucket_chunks_16 [0:63];
    reg [14:0] cnt_bucket_chunks_17 [0:63];
    reg [14:0] cnt_bucket_chunks_18 [0:63];
    reg [14:0] cnt_bucket_chunks_19 [0:63];
    reg [14:0] cnt_bucket_chunks_20 [0:63];
    reg [14:0] cnt_bucket_chunks_21 [0:63];
    reg [14:0] cnt_bucket_chunks_22 [0:63];
    reg [14:0] cnt_bucket_chunks_23 [0:63];
    reg [14:0] cnt_bucket_chunks_24 [0:63];
    reg [14:0] cnt_bucket_chunks_25 [0:63];
    reg [14:0] cnt_bucket_chunks_26 [0:63];
    reg [14:0] cnt_bucket_chunks_27 [0:63];
    reg [14:0] cnt_bucket_chunks_28 [0:63];
    reg [14:0] cnt_bucket_chunks_29 [0:63];
    reg [14:0] cnt_bucket_chunks_30 [0:63];
    reg [14:0] cnt_bucket_chunks_31 [0:63];
    reg [14:0] cnt_bucket_chunks_32 [0:63];
    reg [14:0] cnt_bucket_chunks_33 [0:63];
    reg [14:0] cnt_bucket_chunks_34 [0:63];
    reg [14:0] cnt_bucket_chunks_35 [0:63];
    reg [14:0] cnt_bucket_chunks_36 [0:63];
    reg [14:0] cnt_bucket_chunks_37 [0:63];
    reg [14:0] cnt_bucket_chunks_38 [0:63];
    reg [14:0] cnt_bucket_chunks_39 [0:63];
    reg [14:0] cnt_bucket_chunks_40 [0:63];
    reg [14:0] cnt_bucket_chunks_41 [0:63];
    reg [14:0] cnt_bucket_chunks_42 [0:63];

    wire cnt_bucket_chunks_0_we0, cnt_bucket_chunks_0_we1;
    wire [5:0] cnt_bucket_chunks_0_address0, cnt_bucket_chunks_0_address1;
    wire [14:0] cnt_bucket_chunks_0_d0, cnt_bucket_chunks_0_d1;
    reg [14:0] cnt_bucket_chunks_0_q0, cnt_bucket_chunks_0_q1;
    
    wire cnt_bucket_chunks_1_we0, cnt_bucket_chunks_1_we1;
    wire [5:0] cnt_bucket_chunks_1_address0, cnt_bucket_chunks_1_address1;
    wire [14:0] cnt_bucket_chunks_1_d0, cnt_bucket_chunks_1_d1;
    reg [14:0] cnt_bucket_chunks_1_q0, cnt_bucket_chunks_1_q1;
    
    wire cnt_bucket_chunks_2_we0, cnt_bucket_chunks_2_we1;
    wire [5:0] cnt_bucket_chunks_2_address0, cnt_bucket_chunks_2_address1;
    wire [14:0] cnt_bucket_chunks_2_d0, cnt_bucket_chunks_2_d1;
    reg [14:0] cnt_bucket_chunks_2_q0, cnt_bucket_chunks_2_q1;
    
    wire cnt_bucket_chunks_3_we0, cnt_bucket_chunks_3_we1;
    wire [5:0] cnt_bucket_chunks_3_address0, cnt_bucket_chunks_3_address1;
    wire [14:0] cnt_bucket_chunks_3_d0, cnt_bucket_chunks_3_d1;
    reg [14:0] cnt_bucket_chunks_3_q0, cnt_bucket_chunks_3_q1;
    
    wire cnt_bucket_chunks_4_we0, cnt_bucket_chunks_4_we1;
    wire [5:0] cnt_bucket_chunks_4_address0, cnt_bucket_chunks_4_address1;
    wire [14:0] cnt_bucket_chunks_4_d0, cnt_bucket_chunks_4_d1;
    reg [14:0] cnt_bucket_chunks_4_q0, cnt_bucket_chunks_4_q1;
    
    wire cnt_bucket_chunks_5_we0, cnt_bucket_chunks_5_we1;
    wire [5:0] cnt_bucket_chunks_5_address0, cnt_bucket_chunks_5_address1;
    wire [14:0] cnt_bucket_chunks_5_d0, cnt_bucket_chunks_5_d1;
    reg [14:0] cnt_bucket_chunks_5_q0, cnt_bucket_chunks_5_q1;
    
    wire cnt_bucket_chunks_6_we0, cnt_bucket_chunks_6_we1;
    wire [5:0] cnt_bucket_chunks_6_address0, cnt_bucket_chunks_6_address1;
    wire [14:0] cnt_bucket_chunks_6_d0, cnt_bucket_chunks_6_d1;
    reg [14:0] cnt_bucket_chunks_6_q0, cnt_bucket_chunks_6_q1;
    
    wire cnt_bucket_chunks_7_we0, cnt_bucket_chunks_7_we1;
    wire [5:0] cnt_bucket_chunks_7_address0, cnt_bucket_chunks_7_address1;
    wire [14:0] cnt_bucket_chunks_7_d0, cnt_bucket_chunks_7_d1;
    reg [14:0] cnt_bucket_chunks_7_q0, cnt_bucket_chunks_7_q1;
    
    wire cnt_bucket_chunks_8_we0, cnt_bucket_chunks_8_we1;
    wire [5:0] cnt_bucket_chunks_8_address0, cnt_bucket_chunks_8_address1;
    wire [14:0] cnt_bucket_chunks_8_d0, cnt_bucket_chunks_8_d1;
    reg [14:0] cnt_bucket_chunks_8_q0, cnt_bucket_chunks_8_q1;
    
    wire cnt_bucket_chunks_9_we0, cnt_bucket_chunks_9_we1;
    wire [5:0] cnt_bucket_chunks_9_address0, cnt_bucket_chunks_9_address1;
    wire [14:0] cnt_bucket_chunks_9_d0, cnt_bucket_chunks_9_d1;
    reg [14:0] cnt_bucket_chunks_9_q0, cnt_bucket_chunks_9_q1;
    
    wire cnt_bucket_chunks_10_we0, cnt_bucket_chunks_10_we1;
    wire [5:0] cnt_bucket_chunks_10_address0, cnt_bucket_chunks_10_address1;
    wire [14:0] cnt_bucket_chunks_10_d0, cnt_bucket_chunks_10_d1;
    reg [14:0] cnt_bucket_chunks_10_q0, cnt_bucket_chunks_10_q1;
    
    wire cnt_bucket_chunks_11_we0, cnt_bucket_chunks_11_we1;
    wire [5:0] cnt_bucket_chunks_11_address0, cnt_bucket_chunks_11_address1;
    wire [14:0] cnt_bucket_chunks_11_d0, cnt_bucket_chunks_11_d1;
    reg [14:0] cnt_bucket_chunks_11_q0, cnt_bucket_chunks_11_q1;
    
    wire cnt_bucket_chunks_12_we0, cnt_bucket_chunks_12_we1;
    wire [5:0] cnt_bucket_chunks_12_address0, cnt_bucket_chunks_12_address1;
    wire [14:0] cnt_bucket_chunks_12_d0, cnt_bucket_chunks_12_d1;
    reg [14:0] cnt_bucket_chunks_12_q0, cnt_bucket_chunks_12_q1;
    
    wire cnt_bucket_chunks_13_we0, cnt_bucket_chunks_13_we1;
    wire [5:0] cnt_bucket_chunks_13_address0, cnt_bucket_chunks_13_address1;
    wire [14:0] cnt_bucket_chunks_13_d0, cnt_bucket_chunks_13_d1;
    reg [14:0] cnt_bucket_chunks_13_q0, cnt_bucket_chunks_13_q1;
    
    wire cnt_bucket_chunks_14_we0, cnt_bucket_chunks_14_we1;
    wire [5:0] cnt_bucket_chunks_14_address0, cnt_bucket_chunks_14_address1;
    wire [14:0] cnt_bucket_chunks_14_d0, cnt_bucket_chunks_14_d1;
    reg [14:0] cnt_bucket_chunks_14_q0, cnt_bucket_chunks_14_q1;
    
    wire cnt_bucket_chunks_15_we0, cnt_bucket_chunks_15_we1;
    wire [5:0] cnt_bucket_chunks_15_address0, cnt_bucket_chunks_15_address1;
    wire [14:0] cnt_bucket_chunks_15_d0, cnt_bucket_chunks_15_d1;
    reg [14:0] cnt_bucket_chunks_15_q0, cnt_bucket_chunks_15_q1;
    
    wire cnt_bucket_chunks_16_we0, cnt_bucket_chunks_16_we1;
    wire [5:0] cnt_bucket_chunks_16_address0, cnt_bucket_chunks_16_address1;
    wire [14:0] cnt_bucket_chunks_16_d0, cnt_bucket_chunks_16_d1;
    reg [14:0] cnt_bucket_chunks_16_q0, cnt_bucket_chunks_16_q1;
    
    wire cnt_bucket_chunks_17_we0, cnt_bucket_chunks_17_we1;
    wire [5:0] cnt_bucket_chunks_17_address0, cnt_bucket_chunks_17_address1;
    wire [14:0] cnt_bucket_chunks_17_d0, cnt_bucket_chunks_17_d1;
    reg [14:0] cnt_bucket_chunks_17_q0, cnt_bucket_chunks_17_q1;
    
    wire cnt_bucket_chunks_18_we0, cnt_bucket_chunks_18_we1;
    wire [5:0] cnt_bucket_chunks_18_address0, cnt_bucket_chunks_18_address1;
    wire [14:0] cnt_bucket_chunks_18_d0, cnt_bucket_chunks_18_d1;
    reg [14:0] cnt_bucket_chunks_18_q0, cnt_bucket_chunks_18_q1;
    
    wire cnt_bucket_chunks_19_we0, cnt_bucket_chunks_19_we1;
    wire [5:0] cnt_bucket_chunks_19_address0, cnt_bucket_chunks_19_address1;
    wire [14:0] cnt_bucket_chunks_19_d0, cnt_bucket_chunks_19_d1;
    reg [14:0] cnt_bucket_chunks_19_q0, cnt_bucket_chunks_19_q1;
    
    wire cnt_bucket_chunks_20_we0, cnt_bucket_chunks_20_we1;
    wire [5:0] cnt_bucket_chunks_20_address0, cnt_bucket_chunks_20_address1;
    wire [14:0] cnt_bucket_chunks_20_d0, cnt_bucket_chunks_20_d1;
    reg [14:0] cnt_bucket_chunks_20_q0, cnt_bucket_chunks_20_q1;
    
    wire cnt_bucket_chunks_21_we0, cnt_bucket_chunks_21_we1;
    wire [5:0] cnt_bucket_chunks_21_address0, cnt_bucket_chunks_21_address1;
    wire [14:0] cnt_bucket_chunks_21_d0, cnt_bucket_chunks_21_d1;
    reg [14:0] cnt_bucket_chunks_21_q0, cnt_bucket_chunks_21_q1;
    
    wire cnt_bucket_chunks_22_we0, cnt_bucket_chunks_22_we1;
    wire [5:0] cnt_bucket_chunks_22_address0, cnt_bucket_chunks_22_address1;
    wire [14:0] cnt_bucket_chunks_22_d0, cnt_bucket_chunks_22_d1;
    reg [14:0] cnt_bucket_chunks_22_q0, cnt_bucket_chunks_22_q1;
    
    wire cnt_bucket_chunks_23_we0, cnt_bucket_chunks_23_we1;
    wire [5:0] cnt_bucket_chunks_23_address0, cnt_bucket_chunks_23_address1;
    wire [14:0] cnt_bucket_chunks_23_d0, cnt_bucket_chunks_23_d1;
    reg [14:0] cnt_bucket_chunks_23_q0, cnt_bucket_chunks_23_q1;
    
    wire cnt_bucket_chunks_24_we0, cnt_bucket_chunks_24_we1;
    wire [5:0] cnt_bucket_chunks_24_address0, cnt_bucket_chunks_24_address1;
    wire [14:0] cnt_bucket_chunks_24_d0, cnt_bucket_chunks_24_d1;
    reg [14:0] cnt_bucket_chunks_24_q0, cnt_bucket_chunks_24_q1;
    
    wire cnt_bucket_chunks_25_we0, cnt_bucket_chunks_25_we1;
    wire [5:0] cnt_bucket_chunks_25_address0, cnt_bucket_chunks_25_address1;
    wire [14:0] cnt_bucket_chunks_25_d0, cnt_bucket_chunks_25_d1;
    reg [14:0] cnt_bucket_chunks_25_q0, cnt_bucket_chunks_25_q1;
    
    wire cnt_bucket_chunks_26_we0, cnt_bucket_chunks_26_we1;
    wire [5:0] cnt_bucket_chunks_26_address0, cnt_bucket_chunks_26_address1;
    wire [14:0] cnt_bucket_chunks_26_d0, cnt_bucket_chunks_26_d1;
    reg [14:0] cnt_bucket_chunks_26_q0, cnt_bucket_chunks_26_q1;
    
    wire cnt_bucket_chunks_27_we0, cnt_bucket_chunks_27_we1;
    wire [5:0] cnt_bucket_chunks_27_address0, cnt_bucket_chunks_27_address1;
    wire [14:0] cnt_bucket_chunks_27_d0, cnt_bucket_chunks_27_d1;
    reg [14:0] cnt_bucket_chunks_27_q0, cnt_bucket_chunks_27_q1;
    
    wire cnt_bucket_chunks_28_we0, cnt_bucket_chunks_28_we1;
    wire [5:0] cnt_bucket_chunks_28_address0, cnt_bucket_chunks_28_address1;
    wire [14:0] cnt_bucket_chunks_28_d0, cnt_bucket_chunks_28_d1;
    reg [14:0] cnt_bucket_chunks_28_q0, cnt_bucket_chunks_28_q1;
    
    wire cnt_bucket_chunks_29_we0, cnt_bucket_chunks_29_we1;
    wire [5:0] cnt_bucket_chunks_29_address0, cnt_bucket_chunks_29_address1;
    wire [14:0] cnt_bucket_chunks_29_d0, cnt_bucket_chunks_29_d1;
    reg [14:0] cnt_bucket_chunks_29_q0, cnt_bucket_chunks_29_q1;
    
    wire cnt_bucket_chunks_30_we0, cnt_bucket_chunks_30_we1;
    wire [5:0] cnt_bucket_chunks_30_address0, cnt_bucket_chunks_30_address1;
    wire [14:0] cnt_bucket_chunks_30_d0, cnt_bucket_chunks_30_d1;
    reg [14:0] cnt_bucket_chunks_30_q0, cnt_bucket_chunks_30_q1;
    
    wire cnt_bucket_chunks_31_we0, cnt_bucket_chunks_31_we1;
    wire [5:0] cnt_bucket_chunks_31_address0, cnt_bucket_chunks_31_address1;
    wire [14:0] cnt_bucket_chunks_31_d0, cnt_bucket_chunks_31_d1;
    reg [14:0] cnt_bucket_chunks_31_q0, cnt_bucket_chunks_31_q1;
    
    wire cnt_bucket_chunks_32_we0, cnt_bucket_chunks_32_we1;
    wire [5:0] cnt_bucket_chunks_32_address0, cnt_bucket_chunks_32_address1;
    wire [14:0] cnt_bucket_chunks_32_d0, cnt_bucket_chunks_32_d1;
    reg [14:0] cnt_bucket_chunks_32_q0, cnt_bucket_chunks_32_q1;
    
    wire cnt_bucket_chunks_33_we0, cnt_bucket_chunks_33_we1;
    wire [5:0] cnt_bucket_chunks_33_address0, cnt_bucket_chunks_33_address1;
    wire [14:0] cnt_bucket_chunks_33_d0, cnt_bucket_chunks_33_d1;
    reg [14:0] cnt_bucket_chunks_33_q0, cnt_bucket_chunks_33_q1;
    
    wire cnt_bucket_chunks_34_we0, cnt_bucket_chunks_34_we1;
    wire [5:0] cnt_bucket_chunks_34_address0, cnt_bucket_chunks_34_address1;
    wire [14:0] cnt_bucket_chunks_34_d0, cnt_bucket_chunks_34_d1;
    reg [14:0] cnt_bucket_chunks_34_q0, cnt_bucket_chunks_34_q1;
    
    wire cnt_bucket_chunks_35_we0, cnt_bucket_chunks_35_we1;
    wire [5:0] cnt_bucket_chunks_35_address0, cnt_bucket_chunks_35_address1;
    wire [14:0] cnt_bucket_chunks_35_d0, cnt_bucket_chunks_35_d1;
    reg [14:0] cnt_bucket_chunks_35_q0, cnt_bucket_chunks_35_q1;
    
    wire cnt_bucket_chunks_36_we0, cnt_bucket_chunks_36_we1;
    wire [5:0] cnt_bucket_chunks_36_address0, cnt_bucket_chunks_36_address1;
    wire [14:0] cnt_bucket_chunks_36_d0, cnt_bucket_chunks_36_d1;
    reg [14:0] cnt_bucket_chunks_36_q0, cnt_bucket_chunks_36_q1;
    
    wire cnt_bucket_chunks_37_we0, cnt_bucket_chunks_37_we1;
    wire [5:0] cnt_bucket_chunks_37_address0, cnt_bucket_chunks_37_address1;
    wire [14:0] cnt_bucket_chunks_37_d0, cnt_bucket_chunks_37_d1;
    reg [14:0] cnt_bucket_chunks_37_q0, cnt_bucket_chunks_37_q1;
    
    wire cnt_bucket_chunks_38_we0, cnt_bucket_chunks_38_we1;
    wire [5:0] cnt_bucket_chunks_38_address0, cnt_bucket_chunks_38_address1;
    wire [14:0] cnt_bucket_chunks_38_d0, cnt_bucket_chunks_38_d1;
    reg [14:0] cnt_bucket_chunks_38_q0, cnt_bucket_chunks_38_q1;
    
    wire cnt_bucket_chunks_39_we0, cnt_bucket_chunks_39_we1;
    wire [5:0] cnt_bucket_chunks_39_address0, cnt_bucket_chunks_39_address1;
    wire [14:0] cnt_bucket_chunks_39_d0, cnt_bucket_chunks_39_d1;
    reg [14:0] cnt_bucket_chunks_39_q0, cnt_bucket_chunks_39_q1;
    
    wire cnt_bucket_chunks_40_we0, cnt_bucket_chunks_40_we1;
    wire [5:0] cnt_bucket_chunks_40_address0, cnt_bucket_chunks_40_address1;
    wire [14:0] cnt_bucket_chunks_40_d0, cnt_bucket_chunks_40_d1;
    reg [14:0] cnt_bucket_chunks_40_q0, cnt_bucket_chunks_40_q1;
    
    wire cnt_bucket_chunks_41_we0, cnt_bucket_chunks_41_we1;
    wire [5:0] cnt_bucket_chunks_41_address0, cnt_bucket_chunks_41_address1;
    wire [14:0] cnt_bucket_chunks_41_d0, cnt_bucket_chunks_41_d1;
    reg [14:0] cnt_bucket_chunks_41_q0, cnt_bucket_chunks_41_q1;
    
    wire cnt_bucket_chunks_42_we0, cnt_bucket_chunks_42_we1;
    wire [5:0] cnt_bucket_chunks_42_address0, cnt_bucket_chunks_42_address1;
    wire [14:0] cnt_bucket_chunks_42_d0, cnt_bucket_chunks_42_d1;
    reg [14:0] cnt_bucket_chunks_42_q0, cnt_bucket_chunks_42_q1;
    

    wire   num_padd_ops_stream_empty_n;
    wire   num_padd_ops_stream_read;
    reg [9:0] read_num_padd_ops;
    wire [14:0] num_padd_ops_test_mem_data;

    wire  [4:0] B_i_address0;
    wire   B_i_ce0;
    wire  [31:0] B_i_d0;
    wire  [31:0] B_i_q0;
    wire   B_i_we0;
    wire  [4:0] B_i_address1;
    wire   B_i_ce1;
    wire  [31:0] B_i_d1;
    wire  [31:0] B_i_q1;
    wire   B_i_we1;

    wire [1535:0] msm_return;
        
    initial begin
        $readmemh("/home/sid/Documents/zprize/msm_cloud_sync/hls_zprize_msm/tester/testcase_8/count_chunk_1",cnt_bucket_chunks_0);
        $readmemh("/home/sid/Documents/zprize/msm_cloud_sync/hls_zprize_msm/tester/testcase_8/count_chunk_2",cnt_bucket_chunks_1);
        $readmemh("/home/sid/Documents/zprize/msm_cloud_sync/hls_zprize_msm/tester/testcase_8/count_chunk_3",cnt_bucket_chunks_2);
        $readmemh("/home/sid/Documents/zprize/msm_cloud_sync/hls_zprize_msm/tester/testcase_8/count_chunk_4",cnt_bucket_chunks_3);
        $readmemh("/home/sid/Documents/zprize/msm_cloud_sync/hls_zprize_msm/tester/testcase_8/count_chunk_5",cnt_bucket_chunks_4);
        $readmemh("/home/sid/Documents/zprize/msm_cloud_sync/hls_zprize_msm/tester/testcase_8/count_chunk_6",cnt_bucket_chunks_5);
        $readmemh("/home/sid/Documents/zprize/msm_cloud_sync/hls_zprize_msm/tester/testcase_8/count_chunk_7",cnt_bucket_chunks_6);
        $readmemh("/home/sid/Documents/zprize/msm_cloud_sync/hls_zprize_msm/tester/testcase_8/count_chunk_8",cnt_bucket_chunks_7);
        $readmemh("/home/sid/Documents/zprize/msm_cloud_sync/hls_zprize_msm/tester/testcase_8/count_chunk_9",cnt_bucket_chunks_8);
        $readmemh("/home/sid/Documents/zprize/msm_cloud_sync/hls_zprize_msm/tester/testcase_8/count_chunk_10",cnt_bucket_chunks_9);
        $readmemh("/home/sid/Documents/zprize/msm_cloud_sync/hls_zprize_msm/tester/testcase_8/count_chunk_11",cnt_bucket_chunks_10);
        $readmemh("/home/sid/Documents/zprize/msm_cloud_sync/hls_zprize_msm/tester/testcase_8/count_chunk_12",cnt_bucket_chunks_11);
        $readmemh("/home/sid/Documents/zprize/msm_cloud_sync/hls_zprize_msm/tester/testcase_8/count_chunk_13",cnt_bucket_chunks_12);
        $readmemh("/home/sid/Documents/zprize/msm_cloud_sync/hls_zprize_msm/tester/testcase_8/count_chunk_14",cnt_bucket_chunks_13);
        $readmemh("/home/sid/Documents/zprize/msm_cloud_sync/hls_zprize_msm/tester/testcase_8/count_chunk_15",cnt_bucket_chunks_14);
        $readmemh("/home/sid/Documents/zprize/msm_cloud_sync/hls_zprize_msm/tester/testcase_8/count_chunk_16",cnt_bucket_chunks_15);
        $readmemh("/home/sid/Documents/zprize/msm_cloud_sync/hls_zprize_msm/tester/testcase_8/count_chunk_17",cnt_bucket_chunks_16);
        $readmemh("/home/sid/Documents/zprize/msm_cloud_sync/hls_zprize_msm/tester/testcase_8/count_chunk_18",cnt_bucket_chunks_17);
        $readmemh("/home/sid/Documents/zprize/msm_cloud_sync/hls_zprize_msm/tester/testcase_8/count_chunk_19",cnt_bucket_chunks_18);
        $readmemh("/home/sid/Documents/zprize/msm_cloud_sync/hls_zprize_msm/tester/testcase_8/count_chunk_20",cnt_bucket_chunks_19);
        $readmemh("/home/sid/Documents/zprize/msm_cloud_sync/hls_zprize_msm/tester/testcase_8/count_chunk_21",cnt_bucket_chunks_20);
        $readmemh("/home/sid/Documents/zprize/msm_cloud_sync/hls_zprize_msm/tester/testcase_8/count_chunk_22",cnt_bucket_chunks_21);
        $readmemh("/home/sid/Documents/zprize/msm_cloud_sync/hls_zprize_msm/tester/testcase_8/count_chunk_23",cnt_bucket_chunks_22);
        $readmemh("/home/sid/Documents/zprize/msm_cloud_sync/hls_zprize_msm/tester/testcase_8/count_chunk_24",cnt_bucket_chunks_23);
        $readmemh("/home/sid/Documents/zprize/msm_cloud_sync/hls_zprize_msm/tester/testcase_8/count_chunk_25",cnt_bucket_chunks_24);
        $readmemh("/home/sid/Documents/zprize/msm_cloud_sync/hls_zprize_msm/tester/testcase_8/count_chunk_26",cnt_bucket_chunks_25);
        $readmemh("/home/sid/Documents/zprize/msm_cloud_sync/hls_zprize_msm/tester/testcase_8/count_chunk_27",cnt_bucket_chunks_26);
        $readmemh("/home/sid/Documents/zprize/msm_cloud_sync/hls_zprize_msm/tester/testcase_8/count_chunk_28",cnt_bucket_chunks_27);
        $readmemh("/home/sid/Documents/zprize/msm_cloud_sync/hls_zprize_msm/tester/testcase_8/count_chunk_29",cnt_bucket_chunks_28);
        $readmemh("/home/sid/Documents/zprize/msm_cloud_sync/hls_zprize_msm/tester/testcase_8/count_chunk_30",cnt_bucket_chunks_29);
        $readmemh("/home/sid/Documents/zprize/msm_cloud_sync/hls_zprize_msm/tester/testcase_8/count_chunk_31",cnt_bucket_chunks_30);
        $readmemh("/home/sid/Documents/zprize/msm_cloud_sync/hls_zprize_msm/tester/testcase_8/count_chunk_32",cnt_bucket_chunks_31);
        $readmemh("/home/sid/Documents/zprize/msm_cloud_sync/hls_zprize_msm/tester/testcase_8/count_chunk_33",cnt_bucket_chunks_32);
        $readmemh("/home/sid/Documents/zprize/msm_cloud_sync/hls_zprize_msm/tester/testcase_8/count_chunk_34",cnt_bucket_chunks_33);
        $readmemh("/home/sid/Documents/zprize/msm_cloud_sync/hls_zprize_msm/tester/testcase_8/count_chunk_35",cnt_bucket_chunks_34);
        $readmemh("/home/sid/Documents/zprize/msm_cloud_sync/hls_zprize_msm/tester/testcase_8/count_chunk_36",cnt_bucket_chunks_35);
        $readmemh("/home/sid/Documents/zprize/msm_cloud_sync/hls_zprize_msm/tester/testcase_8/count_chunk_37",cnt_bucket_chunks_36);
        $readmemh("/home/sid/Documents/zprize/msm_cloud_sync/hls_zprize_msm/tester/testcase_8/count_chunk_38",cnt_bucket_chunks_37);
        $readmemh("/home/sid/Documents/zprize/msm_cloud_sync/hls_zprize_msm/tester/testcase_8/count_chunk_39",cnt_bucket_chunks_38);
        $readmemh("/home/sid/Documents/zprize/msm_cloud_sync/hls_zprize_msm/tester/testcase_8/count_chunk_40",cnt_bucket_chunks_39);
        $readmemh("/home/sid/Documents/zprize/msm_cloud_sync/hls_zprize_msm/tester/testcase_8/count_chunk_41",cnt_bucket_chunks_40);
        $readmemh("/home/sid/Documents/zprize/msm_cloud_sync/hls_zprize_msm/tester/testcase_8/count_chunk_42",cnt_bucket_chunks_41);
        $readmemh("/home/sid/Documents/zprize/msm_cloud_sync/hls_zprize_msm/tester/testcase_8/count_chunk_43",cnt_bucket_chunks_42);
        #5;
        ap_clk<=1'b1;
        ap_start<=1'b0;
        ap_rst = 1'b0;
        read_num_padd_ops<=10'b0;
        #20;
        ap_rst = 1'b1; 
        #200;
        ap_rst=1'b0;
        #20;
        ap_start<=1'b1;     
    end
    
    always #(CLK_PERIOD/2) ap_clk <= ~ap_clk;

    always@(posedge ap_clk) begin
        if(ap_done==1'b1) begin
            ap_start<=1'b0;
        end
    end

    assign num_padd_ops_stream_empty_n = ~(read_num_padd_ops==43);

    always@(posedge ap_clk) begin
        if(num_padd_ops_stream_read)
            read_num_padd_ops <= read_num_padd_ops+1'b1;
    end

    always@(posedge ap_clk) begin
    if(cnt_bucket_chunks_0_we0==1'b1)
        cnt_bucket_chunks_0[cnt_bucket_chunks_0_address0] <= cnt_bucket_chunks_0_d0;
    if(cnt_bucket_chunks_0_we1==1'b1)
        cnt_bucket_chunks_0[cnt_bucket_chunks_0_address1] <= cnt_bucket_chunks_0_d1;
    end
    always@(posedge ap_clk) begin
        cnt_bucket_chunks_0_q0 <= cnt_bucket_chunks_0[cnt_bucket_chunks_0_address0];
        cnt_bucket_chunks_0_q1 <= cnt_bucket_chunks_0[cnt_bucket_chunks_0_address1];
    end
    always@(posedge ap_clk) begin
        if(cnt_bucket_chunks_1_we0==1'b1)
            cnt_bucket_chunks_1[cnt_bucket_chunks_1_address0] <= cnt_bucket_chunks_1_d0;
        if(cnt_bucket_chunks_1_we1==1'b1)
            cnt_bucket_chunks_1[cnt_bucket_chunks_1_address1] <= cnt_bucket_chunks_1_d1;
    end
    always@(posedge ap_clk) begin
        cnt_bucket_chunks_1_q0 <= cnt_bucket_chunks_1[cnt_bucket_chunks_1_address0];
        cnt_bucket_chunks_1_q1 <= cnt_bucket_chunks_1[cnt_bucket_chunks_1_address1];
    end
    always@(posedge ap_clk) begin
        if(cnt_bucket_chunks_2_we0==1'b1)
            cnt_bucket_chunks_2[cnt_bucket_chunks_2_address0] <= cnt_bucket_chunks_2_d0;
        if(cnt_bucket_chunks_2_we1==1'b1)
            cnt_bucket_chunks_2[cnt_bucket_chunks_2_address1] <= cnt_bucket_chunks_2_d1;
    end
    always@(posedge ap_clk) begin
        cnt_bucket_chunks_2_q0 <= cnt_bucket_chunks_2[cnt_bucket_chunks_2_address0];
        cnt_bucket_chunks_2_q1 <= cnt_bucket_chunks_2[cnt_bucket_chunks_2_address1];
    end
    always@(posedge ap_clk) begin
        if(cnt_bucket_chunks_3_we0==1'b1)
            cnt_bucket_chunks_3[cnt_bucket_chunks_3_address0] <= cnt_bucket_chunks_3_d0;
        if(cnt_bucket_chunks_3_we1==1'b1)
            cnt_bucket_chunks_3[cnt_bucket_chunks_3_address1] <= cnt_bucket_chunks_3_d1;
    end
    always@(posedge ap_clk) begin
        cnt_bucket_chunks_3_q0 <= cnt_bucket_chunks_3[cnt_bucket_chunks_3_address0];
        cnt_bucket_chunks_3_q1 <= cnt_bucket_chunks_3[cnt_bucket_chunks_3_address1];
    end
    always@(posedge ap_clk) begin
        if(cnt_bucket_chunks_4_we0==1'b1)
            cnt_bucket_chunks_4[cnt_bucket_chunks_4_address0] <= cnt_bucket_chunks_4_d0;
        if(cnt_bucket_chunks_4_we1==1'b1)
            cnt_bucket_chunks_4[cnt_bucket_chunks_4_address1] <= cnt_bucket_chunks_4_d1;
    end
    always@(posedge ap_clk) begin
        cnt_bucket_chunks_4_q0 <= cnt_bucket_chunks_4[cnt_bucket_chunks_4_address0];
        cnt_bucket_chunks_4_q1 <= cnt_bucket_chunks_4[cnt_bucket_chunks_4_address1];
    end
    always@(posedge ap_clk) begin
        if(cnt_bucket_chunks_5_we0==1'b1)
            cnt_bucket_chunks_5[cnt_bucket_chunks_5_address0] <= cnt_bucket_chunks_5_d0;
        if(cnt_bucket_chunks_5_we1==1'b1)
            cnt_bucket_chunks_5[cnt_bucket_chunks_5_address1] <= cnt_bucket_chunks_5_d1;
    end
    always@(posedge ap_clk) begin
        cnt_bucket_chunks_5_q0 <= cnt_bucket_chunks_5[cnt_bucket_chunks_5_address0];
        cnt_bucket_chunks_5_q1 <= cnt_bucket_chunks_5[cnt_bucket_chunks_5_address1];
    end
    always@(posedge ap_clk) begin
        if(cnt_bucket_chunks_6_we0==1'b1)
            cnt_bucket_chunks_6[cnt_bucket_chunks_6_address0] <= cnt_bucket_chunks_6_d0;
        if(cnt_bucket_chunks_6_we1==1'b1)
            cnt_bucket_chunks_6[cnt_bucket_chunks_6_address1] <= cnt_bucket_chunks_6_d1;
    end
    always@(posedge ap_clk) begin
        cnt_bucket_chunks_6_q0 <= cnt_bucket_chunks_6[cnt_bucket_chunks_6_address0];
        cnt_bucket_chunks_6_q1 <= cnt_bucket_chunks_6[cnt_bucket_chunks_6_address1];
    end
    always@(posedge ap_clk) begin
        if(cnt_bucket_chunks_7_we0==1'b1)
            cnt_bucket_chunks_7[cnt_bucket_chunks_7_address0] <= cnt_bucket_chunks_7_d0;
        if(cnt_bucket_chunks_7_we1==1'b1)
            cnt_bucket_chunks_7[cnt_bucket_chunks_7_address1] <= cnt_bucket_chunks_7_d1;
    end
    always@(posedge ap_clk) begin
        cnt_bucket_chunks_7_q0 <= cnt_bucket_chunks_7[cnt_bucket_chunks_7_address0];
        cnt_bucket_chunks_7_q1 <= cnt_bucket_chunks_7[cnt_bucket_chunks_7_address1];
    end
    always@(posedge ap_clk) begin
        if(cnt_bucket_chunks_8_we0==1'b1)
            cnt_bucket_chunks_8[cnt_bucket_chunks_8_address0] <= cnt_bucket_chunks_8_d0;
        if(cnt_bucket_chunks_8_we1==1'b1)
            cnt_bucket_chunks_8[cnt_bucket_chunks_8_address1] <= cnt_bucket_chunks_8_d1;
    end
    always@(posedge ap_clk) begin
        cnt_bucket_chunks_8_q0 <= cnt_bucket_chunks_8[cnt_bucket_chunks_8_address0];
        cnt_bucket_chunks_8_q1 <= cnt_bucket_chunks_8[cnt_bucket_chunks_8_address1];
    end
    always@(posedge ap_clk) begin
        if(cnt_bucket_chunks_9_we0==1'b1)
            cnt_bucket_chunks_9[cnt_bucket_chunks_9_address0] <= cnt_bucket_chunks_9_d0;
        if(cnt_bucket_chunks_9_we1==1'b1)
            cnt_bucket_chunks_9[cnt_bucket_chunks_9_address1] <= cnt_bucket_chunks_9_d1;
    end
    always@(posedge ap_clk) begin
        cnt_bucket_chunks_9_q0 <= cnt_bucket_chunks_9[cnt_bucket_chunks_9_address0];
        cnt_bucket_chunks_9_q1 <= cnt_bucket_chunks_9[cnt_bucket_chunks_9_address1];
    end
    always@(posedge ap_clk) begin
        if(cnt_bucket_chunks_10_we0==1'b1)
            cnt_bucket_chunks_10[cnt_bucket_chunks_10_address0] <= cnt_bucket_chunks_10_d0;
        if(cnt_bucket_chunks_10_we1==1'b1)
            cnt_bucket_chunks_10[cnt_bucket_chunks_10_address1] <= cnt_bucket_chunks_10_d1;
    end
    always@(posedge ap_clk) begin
        cnt_bucket_chunks_10_q0 <= cnt_bucket_chunks_10[cnt_bucket_chunks_10_address0];
        cnt_bucket_chunks_10_q1 <= cnt_bucket_chunks_10[cnt_bucket_chunks_10_address1];
    end
    always@(posedge ap_clk) begin
        if(cnt_bucket_chunks_11_we0==1'b1)
            cnt_bucket_chunks_11[cnt_bucket_chunks_11_address0] <= cnt_bucket_chunks_11_d0;
        if(cnt_bucket_chunks_11_we1==1'b1)
            cnt_bucket_chunks_11[cnt_bucket_chunks_11_address1] <= cnt_bucket_chunks_11_d1;
    end
    always@(posedge ap_clk) begin
        cnt_bucket_chunks_11_q0 <= cnt_bucket_chunks_11[cnt_bucket_chunks_11_address0];
        cnt_bucket_chunks_11_q1 <= cnt_bucket_chunks_11[cnt_bucket_chunks_11_address1];
    end
    always@(posedge ap_clk) begin
        if(cnt_bucket_chunks_12_we0==1'b1)
            cnt_bucket_chunks_12[cnt_bucket_chunks_12_address0] <= cnt_bucket_chunks_12_d0;
        if(cnt_bucket_chunks_12_we1==1'b1)
            cnt_bucket_chunks_12[cnt_bucket_chunks_12_address1] <= cnt_bucket_chunks_12_d1;
    end
    always@(posedge ap_clk) begin
        cnt_bucket_chunks_12_q0 <= cnt_bucket_chunks_12[cnt_bucket_chunks_12_address0];
        cnt_bucket_chunks_12_q1 <= cnt_bucket_chunks_12[cnt_bucket_chunks_12_address1];
    end
    always@(posedge ap_clk) begin
        if(cnt_bucket_chunks_13_we0==1'b1)
            cnt_bucket_chunks_13[cnt_bucket_chunks_13_address0] <= cnt_bucket_chunks_13_d0;
        if(cnt_bucket_chunks_13_we1==1'b1)
            cnt_bucket_chunks_13[cnt_bucket_chunks_13_address1] <= cnt_bucket_chunks_13_d1;
    end
    always@(posedge ap_clk) begin
        cnt_bucket_chunks_13_q0 <= cnt_bucket_chunks_13[cnt_bucket_chunks_13_address0];
        cnt_bucket_chunks_13_q1 <= cnt_bucket_chunks_13[cnt_bucket_chunks_13_address1];
    end
    always@(posedge ap_clk) begin
        if(cnt_bucket_chunks_14_we0==1'b1)
            cnt_bucket_chunks_14[cnt_bucket_chunks_14_address0] <= cnt_bucket_chunks_14_d0;
        if(cnt_bucket_chunks_14_we1==1'b1)
            cnt_bucket_chunks_14[cnt_bucket_chunks_14_address1] <= cnt_bucket_chunks_14_d1;
    end
    always@(posedge ap_clk) begin
        cnt_bucket_chunks_14_q0 <= cnt_bucket_chunks_14[cnt_bucket_chunks_14_address0];
        cnt_bucket_chunks_14_q1 <= cnt_bucket_chunks_14[cnt_bucket_chunks_14_address1];
    end
    always@(posedge ap_clk) begin
        if(cnt_bucket_chunks_15_we0==1'b1)
            cnt_bucket_chunks_15[cnt_bucket_chunks_15_address0] <= cnt_bucket_chunks_15_d0;
        if(cnt_bucket_chunks_15_we1==1'b1)
            cnt_bucket_chunks_15[cnt_bucket_chunks_15_address1] <= cnt_bucket_chunks_15_d1;
    end
    always@(posedge ap_clk) begin
        cnt_bucket_chunks_15_q0 <= cnt_bucket_chunks_15[cnt_bucket_chunks_15_address0];
        cnt_bucket_chunks_15_q1 <= cnt_bucket_chunks_15[cnt_bucket_chunks_15_address1];
    end
    always@(posedge ap_clk) begin
        if(cnt_bucket_chunks_16_we0==1'b1)
            cnt_bucket_chunks_16[cnt_bucket_chunks_16_address0] <= cnt_bucket_chunks_16_d0;
        if(cnt_bucket_chunks_16_we1==1'b1)
            cnt_bucket_chunks_16[cnt_bucket_chunks_16_address1] <= cnt_bucket_chunks_16_d1;
    end
    always@(posedge ap_clk) begin
        cnt_bucket_chunks_16_q0 <= cnt_bucket_chunks_16[cnt_bucket_chunks_16_address0];
        cnt_bucket_chunks_16_q1 <= cnt_bucket_chunks_16[cnt_bucket_chunks_16_address1];
    end
    always@(posedge ap_clk) begin
        if(cnt_bucket_chunks_17_we0==1'b1)
            cnt_bucket_chunks_17[cnt_bucket_chunks_17_address0] <= cnt_bucket_chunks_17_d0;
        if(cnt_bucket_chunks_17_we1==1'b1)
            cnt_bucket_chunks_17[cnt_bucket_chunks_17_address1] <= cnt_bucket_chunks_17_d1;
    end
    always@(posedge ap_clk) begin
        cnt_bucket_chunks_17_q0 <= cnt_bucket_chunks_17[cnt_bucket_chunks_17_address0];
        cnt_bucket_chunks_17_q1 <= cnt_bucket_chunks_17[cnt_bucket_chunks_17_address1];
    end
    always@(posedge ap_clk) begin
        if(cnt_bucket_chunks_18_we0==1'b1)
            cnt_bucket_chunks_18[cnt_bucket_chunks_18_address0] <= cnt_bucket_chunks_18_d0;
        if(cnt_bucket_chunks_18_we1==1'b1)
            cnt_bucket_chunks_18[cnt_bucket_chunks_18_address1] <= cnt_bucket_chunks_18_d1;
    end
    always@(posedge ap_clk) begin
        cnt_bucket_chunks_18_q0 <= cnt_bucket_chunks_18[cnt_bucket_chunks_18_address0];
        cnt_bucket_chunks_18_q1 <= cnt_bucket_chunks_18[cnt_bucket_chunks_18_address1];
    end
    always@(posedge ap_clk) begin
        if(cnt_bucket_chunks_19_we0==1'b1)
            cnt_bucket_chunks_19[cnt_bucket_chunks_19_address0] <= cnt_bucket_chunks_19_d0;
        if(cnt_bucket_chunks_19_we1==1'b1)
            cnt_bucket_chunks_19[cnt_bucket_chunks_19_address1] <= cnt_bucket_chunks_19_d1;
    end
    always@(posedge ap_clk) begin
        cnt_bucket_chunks_19_q0 <= cnt_bucket_chunks_19[cnt_bucket_chunks_19_address0];
        cnt_bucket_chunks_19_q1 <= cnt_bucket_chunks_19[cnt_bucket_chunks_19_address1];
    end
    always@(posedge ap_clk) begin
        if(cnt_bucket_chunks_20_we0==1'b1)
            cnt_bucket_chunks_20[cnt_bucket_chunks_20_address0] <= cnt_bucket_chunks_20_d0;
        if(cnt_bucket_chunks_20_we1==1'b1)
            cnt_bucket_chunks_20[cnt_bucket_chunks_20_address1] <= cnt_bucket_chunks_20_d1;
    end
    always@(posedge ap_clk) begin
        cnt_bucket_chunks_20_q0 <= cnt_bucket_chunks_20[cnt_bucket_chunks_20_address0];
        cnt_bucket_chunks_20_q1 <= cnt_bucket_chunks_20[cnt_bucket_chunks_20_address1];
    end
    always@(posedge ap_clk) begin
        if(cnt_bucket_chunks_21_we0==1'b1)
            cnt_bucket_chunks_21[cnt_bucket_chunks_21_address0] <= cnt_bucket_chunks_21_d0;
        if(cnt_bucket_chunks_21_we1==1'b1)
            cnt_bucket_chunks_21[cnt_bucket_chunks_21_address1] <= cnt_bucket_chunks_21_d1;
    end
    always@(posedge ap_clk) begin
        cnt_bucket_chunks_21_q0 <= cnt_bucket_chunks_21[cnt_bucket_chunks_21_address0];
        cnt_bucket_chunks_21_q1 <= cnt_bucket_chunks_21[cnt_bucket_chunks_21_address1];
    end
    always@(posedge ap_clk) begin
        if(cnt_bucket_chunks_22_we0==1'b1)
            cnt_bucket_chunks_22[cnt_bucket_chunks_22_address0] <= cnt_bucket_chunks_22_d0;
        if(cnt_bucket_chunks_22_we1==1'b1)
            cnt_bucket_chunks_22[cnt_bucket_chunks_22_address1] <= cnt_bucket_chunks_22_d1;
    end
    always@(posedge ap_clk) begin
        cnt_bucket_chunks_22_q0 <= cnt_bucket_chunks_22[cnt_bucket_chunks_22_address0];
        cnt_bucket_chunks_22_q1 <= cnt_bucket_chunks_22[cnt_bucket_chunks_22_address1];
    end
    always@(posedge ap_clk) begin
        if(cnt_bucket_chunks_23_we0==1'b1)
            cnt_bucket_chunks_23[cnt_bucket_chunks_23_address0] <= cnt_bucket_chunks_23_d0;
        if(cnt_bucket_chunks_23_we1==1'b1)
            cnt_bucket_chunks_23[cnt_bucket_chunks_23_address1] <= cnt_bucket_chunks_23_d1;
    end
    always@(posedge ap_clk) begin
        cnt_bucket_chunks_23_q0 <= cnt_bucket_chunks_23[cnt_bucket_chunks_23_address0];
        cnt_bucket_chunks_23_q1 <= cnt_bucket_chunks_23[cnt_bucket_chunks_23_address1];
    end
    always@(posedge ap_clk) begin
        if(cnt_bucket_chunks_24_we0==1'b1)
            cnt_bucket_chunks_24[cnt_bucket_chunks_24_address0] <= cnt_bucket_chunks_24_d0;
        if(cnt_bucket_chunks_24_we1==1'b1)
            cnt_bucket_chunks_24[cnt_bucket_chunks_24_address1] <= cnt_bucket_chunks_24_d1;
    end
    always@(posedge ap_clk) begin
        cnt_bucket_chunks_24_q0 <= cnt_bucket_chunks_24[cnt_bucket_chunks_24_address0];
        cnt_bucket_chunks_24_q1 <= cnt_bucket_chunks_24[cnt_bucket_chunks_24_address1];
    end
    always@(posedge ap_clk) begin
        if(cnt_bucket_chunks_25_we0==1'b1)
            cnt_bucket_chunks_25[cnt_bucket_chunks_25_address0] <= cnt_bucket_chunks_25_d0;
        if(cnt_bucket_chunks_25_we1==1'b1)
            cnt_bucket_chunks_25[cnt_bucket_chunks_25_address1] <= cnt_bucket_chunks_25_d1;
    end
    always@(posedge ap_clk) begin
        cnt_bucket_chunks_25_q0 <= cnt_bucket_chunks_25[cnt_bucket_chunks_25_address0];
        cnt_bucket_chunks_25_q1 <= cnt_bucket_chunks_25[cnt_bucket_chunks_25_address1];
    end
    always@(posedge ap_clk) begin
        if(cnt_bucket_chunks_26_we0==1'b1)
            cnt_bucket_chunks_26[cnt_bucket_chunks_26_address0] <= cnt_bucket_chunks_26_d0;
        if(cnt_bucket_chunks_26_we1==1'b1)
            cnt_bucket_chunks_26[cnt_bucket_chunks_26_address1] <= cnt_bucket_chunks_26_d1;
    end
    always@(posedge ap_clk) begin
        cnt_bucket_chunks_26_q0 <= cnt_bucket_chunks_26[cnt_bucket_chunks_26_address0];
        cnt_bucket_chunks_26_q1 <= cnt_bucket_chunks_26[cnt_bucket_chunks_26_address1];
    end
    always@(posedge ap_clk) begin
        if(cnt_bucket_chunks_27_we0==1'b1)
            cnt_bucket_chunks_27[cnt_bucket_chunks_27_address0] <= cnt_bucket_chunks_27_d0;
        if(cnt_bucket_chunks_27_we1==1'b1)
            cnt_bucket_chunks_27[cnt_bucket_chunks_27_address1] <= cnt_bucket_chunks_27_d1;
    end
    always@(posedge ap_clk) begin
        cnt_bucket_chunks_27_q0 <= cnt_bucket_chunks_27[cnt_bucket_chunks_27_address0];
        cnt_bucket_chunks_27_q1 <= cnt_bucket_chunks_27[cnt_bucket_chunks_27_address1];
    end
    always@(posedge ap_clk) begin
        if(cnt_bucket_chunks_28_we0==1'b1)
            cnt_bucket_chunks_28[cnt_bucket_chunks_28_address0] <= cnt_bucket_chunks_28_d0;
        if(cnt_bucket_chunks_28_we1==1'b1)
            cnt_bucket_chunks_28[cnt_bucket_chunks_28_address1] <= cnt_bucket_chunks_28_d1;
    end
    always@(posedge ap_clk) begin
        cnt_bucket_chunks_28_q0 <= cnt_bucket_chunks_28[cnt_bucket_chunks_28_address0];
        cnt_bucket_chunks_28_q1 <= cnt_bucket_chunks_28[cnt_bucket_chunks_28_address1];
    end
    always@(posedge ap_clk) begin
        if(cnt_bucket_chunks_29_we0==1'b1)
            cnt_bucket_chunks_29[cnt_bucket_chunks_29_address0] <= cnt_bucket_chunks_29_d0;
        if(cnt_bucket_chunks_29_we1==1'b1)
            cnt_bucket_chunks_29[cnt_bucket_chunks_29_address1] <= cnt_bucket_chunks_29_d1;
    end
    always@(posedge ap_clk) begin
        cnt_bucket_chunks_29_q0 <= cnt_bucket_chunks_29[cnt_bucket_chunks_29_address0];
        cnt_bucket_chunks_29_q1 <= cnt_bucket_chunks_29[cnt_bucket_chunks_29_address1];
    end
    always@(posedge ap_clk) begin
        if(cnt_bucket_chunks_30_we0==1'b1)
            cnt_bucket_chunks_30[cnt_bucket_chunks_30_address0] <= cnt_bucket_chunks_30_d0;
        if(cnt_bucket_chunks_30_we1==1'b1)
            cnt_bucket_chunks_30[cnt_bucket_chunks_30_address1] <= cnt_bucket_chunks_30_d1;
    end
    always@(posedge ap_clk) begin
        cnt_bucket_chunks_30_q0 <= cnt_bucket_chunks_30[cnt_bucket_chunks_30_address0];
        cnt_bucket_chunks_30_q1 <= cnt_bucket_chunks_30[cnt_bucket_chunks_30_address1];
    end
    always@(posedge ap_clk) begin
        if(cnt_bucket_chunks_31_we0==1'b1)
            cnt_bucket_chunks_31[cnt_bucket_chunks_31_address0] <= cnt_bucket_chunks_31_d0;
        if(cnt_bucket_chunks_31_we1==1'b1)
            cnt_bucket_chunks_31[cnt_bucket_chunks_31_address1] <= cnt_bucket_chunks_31_d1;
    end
    always@(posedge ap_clk) begin
        cnt_bucket_chunks_31_q0 <= cnt_bucket_chunks_31[cnt_bucket_chunks_31_address0];
        cnt_bucket_chunks_31_q1 <= cnt_bucket_chunks_31[cnt_bucket_chunks_31_address1];
    end
    always@(posedge ap_clk) begin
        if(cnt_bucket_chunks_32_we0==1'b1)
            cnt_bucket_chunks_32[cnt_bucket_chunks_32_address0] <= cnt_bucket_chunks_32_d0;
        if(cnt_bucket_chunks_32_we1==1'b1)
            cnt_bucket_chunks_32[cnt_bucket_chunks_32_address1] <= cnt_bucket_chunks_32_d1;
    end
    always@(posedge ap_clk) begin
        cnt_bucket_chunks_32_q0 <= cnt_bucket_chunks_32[cnt_bucket_chunks_32_address0];
        cnt_bucket_chunks_32_q1 <= cnt_bucket_chunks_32[cnt_bucket_chunks_32_address1];
    end
    always@(posedge ap_clk) begin
        if(cnt_bucket_chunks_33_we0==1'b1)
            cnt_bucket_chunks_33[cnt_bucket_chunks_33_address0] <= cnt_bucket_chunks_33_d0;
        if(cnt_bucket_chunks_33_we1==1'b1)
            cnt_bucket_chunks_33[cnt_bucket_chunks_33_address1] <= cnt_bucket_chunks_33_d1;
    end
    always@(posedge ap_clk) begin
        cnt_bucket_chunks_33_q0 <= cnt_bucket_chunks_33[cnt_bucket_chunks_33_address0];
        cnt_bucket_chunks_33_q1 <= cnt_bucket_chunks_33[cnt_bucket_chunks_33_address1];
    end
    always@(posedge ap_clk) begin
        if(cnt_bucket_chunks_34_we0==1'b1)
            cnt_bucket_chunks_34[cnt_bucket_chunks_34_address0] <= cnt_bucket_chunks_34_d0;
        if(cnt_bucket_chunks_34_we1==1'b1)
            cnt_bucket_chunks_34[cnt_bucket_chunks_34_address1] <= cnt_bucket_chunks_34_d1;
    end
    always@(posedge ap_clk) begin
        cnt_bucket_chunks_34_q0 <= cnt_bucket_chunks_34[cnt_bucket_chunks_34_address0];
        cnt_bucket_chunks_34_q1 <= cnt_bucket_chunks_34[cnt_bucket_chunks_34_address1];
    end
    always@(posedge ap_clk) begin
        if(cnt_bucket_chunks_35_we0==1'b1)
            cnt_bucket_chunks_35[cnt_bucket_chunks_35_address0] <= cnt_bucket_chunks_35_d0;
        if(cnt_bucket_chunks_35_we1==1'b1)
            cnt_bucket_chunks_35[cnt_bucket_chunks_35_address1] <= cnt_bucket_chunks_35_d1;
    end
    always@(posedge ap_clk) begin
        cnt_bucket_chunks_35_q0 <= cnt_bucket_chunks_35[cnt_bucket_chunks_35_address0];
        cnt_bucket_chunks_35_q1 <= cnt_bucket_chunks_35[cnt_bucket_chunks_35_address1];
    end
    always@(posedge ap_clk) begin
        if(cnt_bucket_chunks_36_we0==1'b1)
            cnt_bucket_chunks_36[cnt_bucket_chunks_36_address0] <= cnt_bucket_chunks_36_d0;
        if(cnt_bucket_chunks_36_we1==1'b1)
            cnt_bucket_chunks_36[cnt_bucket_chunks_36_address1] <= cnt_bucket_chunks_36_d1;
    end
    always@(posedge ap_clk) begin
        cnt_bucket_chunks_36_q0 <= cnt_bucket_chunks_36[cnt_bucket_chunks_36_address0];
        cnt_bucket_chunks_36_q1 <= cnt_bucket_chunks_36[cnt_bucket_chunks_36_address1];
    end
    always@(posedge ap_clk) begin
        if(cnt_bucket_chunks_37_we0==1'b1)
            cnt_bucket_chunks_37[cnt_bucket_chunks_37_address0] <= cnt_bucket_chunks_37_d0;
        if(cnt_bucket_chunks_37_we1==1'b1)
            cnt_bucket_chunks_37[cnt_bucket_chunks_37_address1] <= cnt_bucket_chunks_37_d1;
    end
    always@(posedge ap_clk) begin
        cnt_bucket_chunks_37_q0 <= cnt_bucket_chunks_37[cnt_bucket_chunks_37_address0];
        cnt_bucket_chunks_37_q1 <= cnt_bucket_chunks_37[cnt_bucket_chunks_37_address1];
    end
    always@(posedge ap_clk) begin
        if(cnt_bucket_chunks_38_we0==1'b1)
            cnt_bucket_chunks_38[cnt_bucket_chunks_38_address0] <= cnt_bucket_chunks_38_d0;
        if(cnt_bucket_chunks_38_we1==1'b1)
            cnt_bucket_chunks_38[cnt_bucket_chunks_38_address1] <= cnt_bucket_chunks_38_d1;
    end
    always@(posedge ap_clk) begin
        cnt_bucket_chunks_38_q0 <= cnt_bucket_chunks_38[cnt_bucket_chunks_38_address0];
        cnt_bucket_chunks_38_q1 <= cnt_bucket_chunks_38[cnt_bucket_chunks_38_address1];
    end
    always@(posedge ap_clk) begin
        if(cnt_bucket_chunks_39_we0==1'b1)
            cnt_bucket_chunks_39[cnt_bucket_chunks_39_address0] <= cnt_bucket_chunks_39_d0;
        if(cnt_bucket_chunks_39_we1==1'b1)
            cnt_bucket_chunks_39[cnt_bucket_chunks_39_address1] <= cnt_bucket_chunks_39_d1;
    end
    always@(posedge ap_clk) begin
        cnt_bucket_chunks_39_q0 <= cnt_bucket_chunks_39[cnt_bucket_chunks_39_address0];
        cnt_bucket_chunks_39_q1 <= cnt_bucket_chunks_39[cnt_bucket_chunks_39_address1];
    end
    always@(posedge ap_clk) begin
        if(cnt_bucket_chunks_40_we0==1'b1)
            cnt_bucket_chunks_40[cnt_bucket_chunks_40_address0] <= cnt_bucket_chunks_40_d0;
        if(cnt_bucket_chunks_40_we1==1'b1)
            cnt_bucket_chunks_40[cnt_bucket_chunks_40_address1] <= cnt_bucket_chunks_40_d1;
    end
    always@(posedge ap_clk) begin
        cnt_bucket_chunks_40_q0 <= cnt_bucket_chunks_40[cnt_bucket_chunks_40_address0];
        cnt_bucket_chunks_40_q1 <= cnt_bucket_chunks_40[cnt_bucket_chunks_40_address1];
    end
    always@(posedge ap_clk) begin
        if(cnt_bucket_chunks_41_we0==1'b1)
            cnt_bucket_chunks_41[cnt_bucket_chunks_41_address0] <= cnt_bucket_chunks_41_d0;
        if(cnt_bucket_chunks_41_we1==1'b1)
            cnt_bucket_chunks_41[cnt_bucket_chunks_41_address1] <= cnt_bucket_chunks_41_d1;
    end
    always@(posedge ap_clk) begin
        cnt_bucket_chunks_41_q0 <= cnt_bucket_chunks_41[cnt_bucket_chunks_41_address0];
        cnt_bucket_chunks_41_q1 <= cnt_bucket_chunks_41[cnt_bucket_chunks_41_address1];
    end
    always@(posedge ap_clk) begin
        if(cnt_bucket_chunks_42_we0==1'b1)
            cnt_bucket_chunks_42[cnt_bucket_chunks_42_address0] <= cnt_bucket_chunks_42_d0;
        if(cnt_bucket_chunks_42_we1==1'b1)
            cnt_bucket_chunks_42[cnt_bucket_chunks_42_address1] <= cnt_bucket_chunks_42_d1;
    end
    always@(posedge ap_clk) begin
        cnt_bucket_chunks_42_q0 <= cnt_bucket_chunks_42[cnt_bucket_chunks_42_address0];
        cnt_bucket_chunks_42_q1 <= cnt_bucket_chunks_42[cnt_bucket_chunks_42_address1];
    end


/* 
ap_local_block, ap_local_deadlock, ap_clk, ap_rst, ap_start, ap_done, ap_idle, ap_ready, P_arr_x_address0, P_arr_x_ce0, P_arr_x_q0, P_arr_y_address0, P_arr_y_ce0, P_arr_y_q0, P_arr_z_address0, P_arr_z_ce0, P_arr_z_q0, K_arr_address0, K_arr_ce0, K_arr_q0, B_i_address0, B_i_ce0, B_i_we0, B_i_d0, B_i_address1, B_i_ce1, B_i_we1, B_i_d1
*/

    top uut(
        .ap_clk(ap_clk),
        .ap_rst(ap_rst),
        .ap_start(ap_start),
        .ap_done(ap_done),
        .ap_idle(ap_idle),
        .ap_ready(ap_ready),
        .P_arr_x_address0(P_arr_x_address0),
        .P_arr_x_ce0(P_arr_x_ce0),
        .P_arr_x_we0(P_arr_x_we0),
        .P_arr_x_q0(P_arr_x_q0),
        .P_arr_x_d0(P_arr_x_d0),
        .P_arr_y_address0(P_arr_y_address0),
        .P_arr_y_ce0(P_arr_y_ce0),
        .P_arr_y_we0(P_arr_y_we0),
        .P_arr_y_q0(P_arr_y_q0),
        .P_arr_y_d0(P_arr_y_d0),
        .P_arr_z_address0(P_arr_z_address0),
        .P_arr_z_ce0(P_arr_z_ce0),
        .P_arr_z_we0(P_arr_z_we0),
        .P_arr_z_q0(P_arr_z_q0),
        .P_arr_z_d0(P_arr_z_d0),
        .P_arr_x_address1(P_arr_x_address1),
        .P_arr_x_ce1(P_arr_x_ce1),
        .P_arr_x_we1(P_arr_x_we1),
        .P_arr_x_q1(P_arr_x_q1),
        .P_arr_x_d1(P_arr_x_d1),
        .P_arr_y_address1(P_arr_y_address1),
        .P_arr_y_ce1(P_arr_y_ce1),
        .P_arr_y_we1(P_arr_y_we1),
        .P_arr_y_q1(P_arr_y_q1),
        .P_arr_y_d1(P_arr_y_d1),
        .P_arr_z_address1(P_arr_z_address1),
        .P_arr_z_ce1(P_arr_z_ce1),
        .P_arr_z_we1(P_arr_z_we1),
        .P_arr_z_q1(P_arr_z_q1),
        .P_arr_z_d1(P_arr_z_d1),
        .K_arr_address0(K_arr_address0),
        .K_arr_ce0(K_arr_ce0),
        .K_arr_we0(K_arr_we0),
        .K_arr_q0(K_arr_q0),
        .K_arr_d0(K_arr_d0),
        // .K_arr_address1(K_arr_address1),
        // .K_arr_ce1(K_arr_ce1),
        // .K_arr_we1(K_arr_we1),
        // .K_arr_q1(K_arr_q1),
        // .K_arr_d1(K_arr_d1),
        .cnt_bucket_chunks_0_address0(cnt_bucket_chunks_0_address0),
        .cnt_bucket_chunks_0_ce0(cnt_bucket_chunks_0_ce0),
        .cnt_bucket_chunks_0_d0(cnt_bucket_chunks_0_d0),
        .cnt_bucket_chunks_0_q0(cnt_bucket_chunks_0_q0),
        .cnt_bucket_chunks_0_we0(cnt_bucket_chunks_0_we0),
        .cnt_bucket_chunks_0_address1(cnt_bucket_chunks_0_address1),
        .cnt_bucket_chunks_0_ce1(cnt_bucket_chunks_0_ce1),
        .cnt_bucket_chunks_0_d1(cnt_bucket_chunks_0_d1),
        .cnt_bucket_chunks_0_q1(cnt_bucket_chunks_0_q1),
        .cnt_bucket_chunks_0_we1(cnt_bucket_chunks_0_we1),
        .cnt_bucket_chunks_1_address0(cnt_bucket_chunks_1_address0),
        .cnt_bucket_chunks_1_ce0(cnt_bucket_chunks_1_ce0),
        .cnt_bucket_chunks_1_d0(cnt_bucket_chunks_1_d0),
        .cnt_bucket_chunks_1_q0(cnt_bucket_chunks_1_q0),
        .cnt_bucket_chunks_1_we0(cnt_bucket_chunks_1_we0),
        .cnt_bucket_chunks_1_address1(cnt_bucket_chunks_1_address1),
        .cnt_bucket_chunks_1_ce1(cnt_bucket_chunks_1_ce1),
        .cnt_bucket_chunks_1_d1(cnt_bucket_chunks_1_d1),
        .cnt_bucket_chunks_1_q1(cnt_bucket_chunks_1_q1),
        .cnt_bucket_chunks_1_we1(cnt_bucket_chunks_1_we1),
        .cnt_bucket_chunks_2_address0(cnt_bucket_chunks_2_address0),
        .cnt_bucket_chunks_2_ce0(cnt_bucket_chunks_2_ce0),
        .cnt_bucket_chunks_2_d0(cnt_bucket_chunks_2_d0),
        .cnt_bucket_chunks_2_q0(cnt_bucket_chunks_2_q0),
        .cnt_bucket_chunks_2_we0(cnt_bucket_chunks_2_we0),
        .cnt_bucket_chunks_2_address1(cnt_bucket_chunks_2_address1),
        .cnt_bucket_chunks_2_ce1(cnt_bucket_chunks_2_ce1),
        .cnt_bucket_chunks_2_d1(cnt_bucket_chunks_2_d1),
        .cnt_bucket_chunks_2_q1(cnt_bucket_chunks_2_q1),
        .cnt_bucket_chunks_2_we1(cnt_bucket_chunks_2_we1),
        .cnt_bucket_chunks_3_address0(cnt_bucket_chunks_3_address0),
        .cnt_bucket_chunks_3_ce0(cnt_bucket_chunks_3_ce0),
        .cnt_bucket_chunks_3_d0(cnt_bucket_chunks_3_d0),
        .cnt_bucket_chunks_3_q0(cnt_bucket_chunks_3_q0),
        .cnt_bucket_chunks_3_we0(cnt_bucket_chunks_3_we0),
        .cnt_bucket_chunks_3_address1(cnt_bucket_chunks_3_address1),
        .cnt_bucket_chunks_3_ce1(cnt_bucket_chunks_3_ce1),
        .cnt_bucket_chunks_3_d1(cnt_bucket_chunks_3_d1),
        .cnt_bucket_chunks_3_q1(cnt_bucket_chunks_3_q1),
        .cnt_bucket_chunks_3_we1(cnt_bucket_chunks_3_we1),
        .cnt_bucket_chunks_4_address0(cnt_bucket_chunks_4_address0),
        .cnt_bucket_chunks_4_ce0(cnt_bucket_chunks_4_ce0),
        .cnt_bucket_chunks_4_d0(cnt_bucket_chunks_4_d0),
        .cnt_bucket_chunks_4_q0(cnt_bucket_chunks_4_q0),
        .cnt_bucket_chunks_4_we0(cnt_bucket_chunks_4_we0),
        .cnt_bucket_chunks_4_address1(cnt_bucket_chunks_4_address1),
        .cnt_bucket_chunks_4_ce1(cnt_bucket_chunks_4_ce1),
        .cnt_bucket_chunks_4_d1(cnt_bucket_chunks_4_d1),
        .cnt_bucket_chunks_4_q1(cnt_bucket_chunks_4_q1),
        .cnt_bucket_chunks_4_we1(cnt_bucket_chunks_4_we1),
        .cnt_bucket_chunks_5_address0(cnt_bucket_chunks_5_address0),
        .cnt_bucket_chunks_5_ce0(cnt_bucket_chunks_5_ce0),
        .cnt_bucket_chunks_5_d0(cnt_bucket_chunks_5_d0),
        .cnt_bucket_chunks_5_q0(cnt_bucket_chunks_5_q0),
        .cnt_bucket_chunks_5_we0(cnt_bucket_chunks_5_we0),
        .cnt_bucket_chunks_5_address1(cnt_bucket_chunks_5_address1),
        .cnt_bucket_chunks_5_ce1(cnt_bucket_chunks_5_ce1),
        .cnt_bucket_chunks_5_d1(cnt_bucket_chunks_5_d1),
        .cnt_bucket_chunks_5_q1(cnt_bucket_chunks_5_q1),
        .cnt_bucket_chunks_5_we1(cnt_bucket_chunks_5_we1),
        .cnt_bucket_chunks_6_address0(cnt_bucket_chunks_6_address0),
        .cnt_bucket_chunks_6_ce0(cnt_bucket_chunks_6_ce0),
        .cnt_bucket_chunks_6_d0(cnt_bucket_chunks_6_d0),
        .cnt_bucket_chunks_6_q0(cnt_bucket_chunks_6_q0),
        .cnt_bucket_chunks_6_we0(cnt_bucket_chunks_6_we0),
        .cnt_bucket_chunks_6_address1(cnt_bucket_chunks_6_address1),
        .cnt_bucket_chunks_6_ce1(cnt_bucket_chunks_6_ce1),
        .cnt_bucket_chunks_6_d1(cnt_bucket_chunks_6_d1),
        .cnt_bucket_chunks_6_q1(cnt_bucket_chunks_6_q1),
        .cnt_bucket_chunks_6_we1(cnt_bucket_chunks_6_we1),
        .cnt_bucket_chunks_7_address0(cnt_bucket_chunks_7_address0),
        .cnt_bucket_chunks_7_ce0(cnt_bucket_chunks_7_ce0),
        .cnt_bucket_chunks_7_d0(cnt_bucket_chunks_7_d0),
        .cnt_bucket_chunks_7_q0(cnt_bucket_chunks_7_q0),
        .cnt_bucket_chunks_7_we0(cnt_bucket_chunks_7_we0),
        .cnt_bucket_chunks_7_address1(cnt_bucket_chunks_7_address1),
        .cnt_bucket_chunks_7_ce1(cnt_bucket_chunks_7_ce1),
        .cnt_bucket_chunks_7_d1(cnt_bucket_chunks_7_d1),
        .cnt_bucket_chunks_7_q1(cnt_bucket_chunks_7_q1),
        .cnt_bucket_chunks_7_we1(cnt_bucket_chunks_7_we1),
        .cnt_bucket_chunks_8_address0(cnt_bucket_chunks_8_address0),
        .cnt_bucket_chunks_8_ce0(cnt_bucket_chunks_8_ce0),
        .cnt_bucket_chunks_8_d0(cnt_bucket_chunks_8_d0),
        .cnt_bucket_chunks_8_q0(cnt_bucket_chunks_8_q0),
        .cnt_bucket_chunks_8_we0(cnt_bucket_chunks_8_we0),
        .cnt_bucket_chunks_8_address1(cnt_bucket_chunks_8_address1),
        .cnt_bucket_chunks_8_ce1(cnt_bucket_chunks_8_ce1),
        .cnt_bucket_chunks_8_d1(cnt_bucket_chunks_8_d1),
        .cnt_bucket_chunks_8_q1(cnt_bucket_chunks_8_q1),
        .cnt_bucket_chunks_8_we1(cnt_bucket_chunks_8_we1),
        .cnt_bucket_chunks_9_address0(cnt_bucket_chunks_9_address0),
        .cnt_bucket_chunks_9_ce0(cnt_bucket_chunks_9_ce0),
        .cnt_bucket_chunks_9_d0(cnt_bucket_chunks_9_d0),
        .cnt_bucket_chunks_9_q0(cnt_bucket_chunks_9_q0),
        .cnt_bucket_chunks_9_we0(cnt_bucket_chunks_9_we0),
        .cnt_bucket_chunks_9_address1(cnt_bucket_chunks_9_address1),
        .cnt_bucket_chunks_9_ce1(cnt_bucket_chunks_9_ce1),
        .cnt_bucket_chunks_9_d1(cnt_bucket_chunks_9_d1),
        .cnt_bucket_chunks_9_q1(cnt_bucket_chunks_9_q1),
        .cnt_bucket_chunks_9_we1(cnt_bucket_chunks_9_we1),
        .cnt_bucket_chunks_10_address0(cnt_bucket_chunks_10_address0),
        .cnt_bucket_chunks_10_ce0(cnt_bucket_chunks_10_ce0),
        .cnt_bucket_chunks_10_d0(cnt_bucket_chunks_10_d0),
        .cnt_bucket_chunks_10_q0(cnt_bucket_chunks_10_q0),
        .cnt_bucket_chunks_10_we0(cnt_bucket_chunks_10_we0),
        .cnt_bucket_chunks_10_address1(cnt_bucket_chunks_10_address1),
        .cnt_bucket_chunks_10_ce1(cnt_bucket_chunks_10_ce1),
        .cnt_bucket_chunks_10_d1(cnt_bucket_chunks_10_d1),
        .cnt_bucket_chunks_10_q1(cnt_bucket_chunks_10_q1),
        .cnt_bucket_chunks_10_we1(cnt_bucket_chunks_10_we1),
        .cnt_bucket_chunks_11_address0(cnt_bucket_chunks_11_address0),
        .cnt_bucket_chunks_11_ce0(cnt_bucket_chunks_11_ce0),
        .cnt_bucket_chunks_11_d0(cnt_bucket_chunks_11_d0),
        .cnt_bucket_chunks_11_q0(cnt_bucket_chunks_11_q0),
        .cnt_bucket_chunks_11_we0(cnt_bucket_chunks_11_we0),
        .cnt_bucket_chunks_11_address1(cnt_bucket_chunks_11_address1),
        .cnt_bucket_chunks_11_ce1(cnt_bucket_chunks_11_ce1),
        .cnt_bucket_chunks_11_d1(cnt_bucket_chunks_11_d1),
        .cnt_bucket_chunks_11_q1(cnt_bucket_chunks_11_q1),
        .cnt_bucket_chunks_11_we1(cnt_bucket_chunks_11_we1),
        .cnt_bucket_chunks_12_address0(cnt_bucket_chunks_12_address0),
        .cnt_bucket_chunks_12_ce0(cnt_bucket_chunks_12_ce0),
        .cnt_bucket_chunks_12_d0(cnt_bucket_chunks_12_d0),
        .cnt_bucket_chunks_12_q0(cnt_bucket_chunks_12_q0),
        .cnt_bucket_chunks_12_we0(cnt_bucket_chunks_12_we0),
        .cnt_bucket_chunks_12_address1(cnt_bucket_chunks_12_address1),
        .cnt_bucket_chunks_12_ce1(cnt_bucket_chunks_12_ce1),
        .cnt_bucket_chunks_12_d1(cnt_bucket_chunks_12_d1),
        .cnt_bucket_chunks_12_q1(cnt_bucket_chunks_12_q1),
        .cnt_bucket_chunks_12_we1(cnt_bucket_chunks_12_we1),
        .cnt_bucket_chunks_13_address0(cnt_bucket_chunks_13_address0),
        .cnt_bucket_chunks_13_ce0(cnt_bucket_chunks_13_ce0),
        .cnt_bucket_chunks_13_d0(cnt_bucket_chunks_13_d0),
        .cnt_bucket_chunks_13_q0(cnt_bucket_chunks_13_q0),
        .cnt_bucket_chunks_13_we0(cnt_bucket_chunks_13_we0),
        .cnt_bucket_chunks_13_address1(cnt_bucket_chunks_13_address1),
        .cnt_bucket_chunks_13_ce1(cnt_bucket_chunks_13_ce1),
        .cnt_bucket_chunks_13_d1(cnt_bucket_chunks_13_d1),
        .cnt_bucket_chunks_13_q1(cnt_bucket_chunks_13_q1),
        .cnt_bucket_chunks_13_we1(cnt_bucket_chunks_13_we1),
        .cnt_bucket_chunks_14_address0(cnt_bucket_chunks_14_address0),
        .cnt_bucket_chunks_14_ce0(cnt_bucket_chunks_14_ce0),
        .cnt_bucket_chunks_14_d0(cnt_bucket_chunks_14_d0),
        .cnt_bucket_chunks_14_q0(cnt_bucket_chunks_14_q0),
        .cnt_bucket_chunks_14_we0(cnt_bucket_chunks_14_we0),
        .cnt_bucket_chunks_14_address1(cnt_bucket_chunks_14_address1),
        .cnt_bucket_chunks_14_ce1(cnt_bucket_chunks_14_ce1),
        .cnt_bucket_chunks_14_d1(cnt_bucket_chunks_14_d1),
        .cnt_bucket_chunks_14_q1(cnt_bucket_chunks_14_q1),
        .cnt_bucket_chunks_14_we1(cnt_bucket_chunks_14_we1),
        .cnt_bucket_chunks_15_address0(cnt_bucket_chunks_15_address0),
        .cnt_bucket_chunks_15_ce0(cnt_bucket_chunks_15_ce0),
        .cnt_bucket_chunks_15_d0(cnt_bucket_chunks_15_d0),
        .cnt_bucket_chunks_15_q0(cnt_bucket_chunks_15_q0),
        .cnt_bucket_chunks_15_we0(cnt_bucket_chunks_15_we0),
        .cnt_bucket_chunks_15_address1(cnt_bucket_chunks_15_address1),
        .cnt_bucket_chunks_15_ce1(cnt_bucket_chunks_15_ce1),
        .cnt_bucket_chunks_15_d1(cnt_bucket_chunks_15_d1),
        .cnt_bucket_chunks_15_q1(cnt_bucket_chunks_15_q1),
        .cnt_bucket_chunks_15_we1(cnt_bucket_chunks_15_we1),
        .cnt_bucket_chunks_16_address0(cnt_bucket_chunks_16_address0),
        .cnt_bucket_chunks_16_ce0(cnt_bucket_chunks_16_ce0),
        .cnt_bucket_chunks_16_d0(cnt_bucket_chunks_16_d0),
        .cnt_bucket_chunks_16_q0(cnt_bucket_chunks_16_q0),
        .cnt_bucket_chunks_16_we0(cnt_bucket_chunks_16_we0),
        .cnt_bucket_chunks_16_address1(cnt_bucket_chunks_16_address1),
        .cnt_bucket_chunks_16_ce1(cnt_bucket_chunks_16_ce1),
        .cnt_bucket_chunks_16_d1(cnt_bucket_chunks_16_d1),
        .cnt_bucket_chunks_16_q1(cnt_bucket_chunks_16_q1),
        .cnt_bucket_chunks_16_we1(cnt_bucket_chunks_16_we1),
        .cnt_bucket_chunks_17_address0(cnt_bucket_chunks_17_address0),
        .cnt_bucket_chunks_17_ce0(cnt_bucket_chunks_17_ce0),
        .cnt_bucket_chunks_17_d0(cnt_bucket_chunks_17_d0),
        .cnt_bucket_chunks_17_q0(cnt_bucket_chunks_17_q0),
        .cnt_bucket_chunks_17_we0(cnt_bucket_chunks_17_we0),
        .cnt_bucket_chunks_17_address1(cnt_bucket_chunks_17_address1),
        .cnt_bucket_chunks_17_ce1(cnt_bucket_chunks_17_ce1),
        .cnt_bucket_chunks_17_d1(cnt_bucket_chunks_17_d1),
        .cnt_bucket_chunks_17_q1(cnt_bucket_chunks_17_q1),
        .cnt_bucket_chunks_17_we1(cnt_bucket_chunks_17_we1),
        .cnt_bucket_chunks_18_address0(cnt_bucket_chunks_18_address0),
        .cnt_bucket_chunks_18_ce0(cnt_bucket_chunks_18_ce0),
        .cnt_bucket_chunks_18_d0(cnt_bucket_chunks_18_d0),
        .cnt_bucket_chunks_18_q0(cnt_bucket_chunks_18_q0),
        .cnt_bucket_chunks_18_we0(cnt_bucket_chunks_18_we0),
        .cnt_bucket_chunks_18_address1(cnt_bucket_chunks_18_address1),
        .cnt_bucket_chunks_18_ce1(cnt_bucket_chunks_18_ce1),
        .cnt_bucket_chunks_18_d1(cnt_bucket_chunks_18_d1),
        .cnt_bucket_chunks_18_q1(cnt_bucket_chunks_18_q1),
        .cnt_bucket_chunks_18_we1(cnt_bucket_chunks_18_we1),
        .cnt_bucket_chunks_19_address0(cnt_bucket_chunks_19_address0),
        .cnt_bucket_chunks_19_ce0(cnt_bucket_chunks_19_ce0),
        .cnt_bucket_chunks_19_d0(cnt_bucket_chunks_19_d0),
        .cnt_bucket_chunks_19_q0(cnt_bucket_chunks_19_q0),
        .cnt_bucket_chunks_19_we0(cnt_bucket_chunks_19_we0),
        .cnt_bucket_chunks_19_address1(cnt_bucket_chunks_19_address1),
        .cnt_bucket_chunks_19_ce1(cnt_bucket_chunks_19_ce1),
        .cnt_bucket_chunks_19_d1(cnt_bucket_chunks_19_d1),
        .cnt_bucket_chunks_19_q1(cnt_bucket_chunks_19_q1),
        .cnt_bucket_chunks_19_we1(cnt_bucket_chunks_19_we1),
        .cnt_bucket_chunks_20_address0(cnt_bucket_chunks_20_address0),
        .cnt_bucket_chunks_20_ce0(cnt_bucket_chunks_20_ce0),
        .cnt_bucket_chunks_20_d0(cnt_bucket_chunks_20_d0),
        .cnt_bucket_chunks_20_q0(cnt_bucket_chunks_20_q0),
        .cnt_bucket_chunks_20_we0(cnt_bucket_chunks_20_we0),
        .cnt_bucket_chunks_20_address1(cnt_bucket_chunks_20_address1),
        .cnt_bucket_chunks_20_ce1(cnt_bucket_chunks_20_ce1),
        .cnt_bucket_chunks_20_d1(cnt_bucket_chunks_20_d1),
        .cnt_bucket_chunks_20_q1(cnt_bucket_chunks_20_q1),
        .cnt_bucket_chunks_20_we1(cnt_bucket_chunks_20_we1),
        .cnt_bucket_chunks_21_address0(cnt_bucket_chunks_21_address0),
        .cnt_bucket_chunks_21_ce0(cnt_bucket_chunks_21_ce0),
        .cnt_bucket_chunks_21_d0(cnt_bucket_chunks_21_d0),
        .cnt_bucket_chunks_21_q0(cnt_bucket_chunks_21_q0),
        .cnt_bucket_chunks_21_we0(cnt_bucket_chunks_21_we0),
        .cnt_bucket_chunks_21_address1(cnt_bucket_chunks_21_address1),
        .cnt_bucket_chunks_21_ce1(cnt_bucket_chunks_21_ce1),
        .cnt_bucket_chunks_21_d1(cnt_bucket_chunks_21_d1),
        .cnt_bucket_chunks_21_q1(cnt_bucket_chunks_21_q1),
        .cnt_bucket_chunks_21_we1(cnt_bucket_chunks_21_we1),
        .cnt_bucket_chunks_22_address0(cnt_bucket_chunks_22_address0),
        .cnt_bucket_chunks_22_ce0(cnt_bucket_chunks_22_ce0),
        .cnt_bucket_chunks_22_d0(cnt_bucket_chunks_22_d0),
        .cnt_bucket_chunks_22_q0(cnt_bucket_chunks_22_q0),
        .cnt_bucket_chunks_22_we0(cnt_bucket_chunks_22_we0),
        .cnt_bucket_chunks_22_address1(cnt_bucket_chunks_22_address1),
        .cnt_bucket_chunks_22_ce1(cnt_bucket_chunks_22_ce1),
        .cnt_bucket_chunks_22_d1(cnt_bucket_chunks_22_d1),
        .cnt_bucket_chunks_22_q1(cnt_bucket_chunks_22_q1),
        .cnt_bucket_chunks_22_we1(cnt_bucket_chunks_22_we1),
        .cnt_bucket_chunks_23_address0(cnt_bucket_chunks_23_address0),
        .cnt_bucket_chunks_23_ce0(cnt_bucket_chunks_23_ce0),
        .cnt_bucket_chunks_23_d0(cnt_bucket_chunks_23_d0),
        .cnt_bucket_chunks_23_q0(cnt_bucket_chunks_23_q0),
        .cnt_bucket_chunks_23_we0(cnt_bucket_chunks_23_we0),
        .cnt_bucket_chunks_23_address1(cnt_bucket_chunks_23_address1),
        .cnt_bucket_chunks_23_ce1(cnt_bucket_chunks_23_ce1),
        .cnt_bucket_chunks_23_d1(cnt_bucket_chunks_23_d1),
        .cnt_bucket_chunks_23_q1(cnt_bucket_chunks_23_q1),
        .cnt_bucket_chunks_23_we1(cnt_bucket_chunks_23_we1),
        .cnt_bucket_chunks_24_address0(cnt_bucket_chunks_24_address0),
        .cnt_bucket_chunks_24_ce0(cnt_bucket_chunks_24_ce0),
        .cnt_bucket_chunks_24_d0(cnt_bucket_chunks_24_d0),
        .cnt_bucket_chunks_24_q0(cnt_bucket_chunks_24_q0),
        .cnt_bucket_chunks_24_we0(cnt_bucket_chunks_24_we0),
        .cnt_bucket_chunks_24_address1(cnt_bucket_chunks_24_address1),
        .cnt_bucket_chunks_24_ce1(cnt_bucket_chunks_24_ce1),
        .cnt_bucket_chunks_24_d1(cnt_bucket_chunks_24_d1),
        .cnt_bucket_chunks_24_q1(cnt_bucket_chunks_24_q1),
        .cnt_bucket_chunks_24_we1(cnt_bucket_chunks_24_we1),
        .cnt_bucket_chunks_25_address0(cnt_bucket_chunks_25_address0),
        .cnt_bucket_chunks_25_ce0(cnt_bucket_chunks_25_ce0),
        .cnt_bucket_chunks_25_d0(cnt_bucket_chunks_25_d0),
        .cnt_bucket_chunks_25_q0(cnt_bucket_chunks_25_q0),
        .cnt_bucket_chunks_25_we0(cnt_bucket_chunks_25_we0),
        .cnt_bucket_chunks_25_address1(cnt_bucket_chunks_25_address1),
        .cnt_bucket_chunks_25_ce1(cnt_bucket_chunks_25_ce1),
        .cnt_bucket_chunks_25_d1(cnt_bucket_chunks_25_d1),
        .cnt_bucket_chunks_25_q1(cnt_bucket_chunks_25_q1),
        .cnt_bucket_chunks_25_we1(cnt_bucket_chunks_25_we1),
        .cnt_bucket_chunks_26_address0(cnt_bucket_chunks_26_address0),
        .cnt_bucket_chunks_26_ce0(cnt_bucket_chunks_26_ce0),
        .cnt_bucket_chunks_26_d0(cnt_bucket_chunks_26_d0),
        .cnt_bucket_chunks_26_q0(cnt_bucket_chunks_26_q0),
        .cnt_bucket_chunks_26_we0(cnt_bucket_chunks_26_we0),
        .cnt_bucket_chunks_26_address1(cnt_bucket_chunks_26_address1),
        .cnt_bucket_chunks_26_ce1(cnt_bucket_chunks_26_ce1),
        .cnt_bucket_chunks_26_d1(cnt_bucket_chunks_26_d1),
        .cnt_bucket_chunks_26_q1(cnt_bucket_chunks_26_q1),
        .cnt_bucket_chunks_26_we1(cnt_bucket_chunks_26_we1),
        .cnt_bucket_chunks_27_address0(cnt_bucket_chunks_27_address0),
        .cnt_bucket_chunks_27_ce0(cnt_bucket_chunks_27_ce0),
        .cnt_bucket_chunks_27_d0(cnt_bucket_chunks_27_d0),
        .cnt_bucket_chunks_27_q0(cnt_bucket_chunks_27_q0),
        .cnt_bucket_chunks_27_we0(cnt_bucket_chunks_27_we0),
        .cnt_bucket_chunks_27_address1(cnt_bucket_chunks_27_address1),
        .cnt_bucket_chunks_27_ce1(cnt_bucket_chunks_27_ce1),
        .cnt_bucket_chunks_27_d1(cnt_bucket_chunks_27_d1),
        .cnt_bucket_chunks_27_q1(cnt_bucket_chunks_27_q1),
        .cnt_bucket_chunks_27_we1(cnt_bucket_chunks_27_we1),
        .cnt_bucket_chunks_28_address0(cnt_bucket_chunks_28_address0),
        .cnt_bucket_chunks_28_ce0(cnt_bucket_chunks_28_ce0),
        .cnt_bucket_chunks_28_d0(cnt_bucket_chunks_28_d0),
        .cnt_bucket_chunks_28_q0(cnt_bucket_chunks_28_q0),
        .cnt_bucket_chunks_28_we0(cnt_bucket_chunks_28_we0),
        .cnt_bucket_chunks_28_address1(cnt_bucket_chunks_28_address1),
        .cnt_bucket_chunks_28_ce1(cnt_bucket_chunks_28_ce1),
        .cnt_bucket_chunks_28_d1(cnt_bucket_chunks_28_d1),
        .cnt_bucket_chunks_28_q1(cnt_bucket_chunks_28_q1),
        .cnt_bucket_chunks_28_we1(cnt_bucket_chunks_28_we1),
        .cnt_bucket_chunks_29_address0(cnt_bucket_chunks_29_address0),
        .cnt_bucket_chunks_29_ce0(cnt_bucket_chunks_29_ce0),
        .cnt_bucket_chunks_29_d0(cnt_bucket_chunks_29_d0),
        .cnt_bucket_chunks_29_q0(cnt_bucket_chunks_29_q0),
        .cnt_bucket_chunks_29_we0(cnt_bucket_chunks_29_we0),
        .cnt_bucket_chunks_29_address1(cnt_bucket_chunks_29_address1),
        .cnt_bucket_chunks_29_ce1(cnt_bucket_chunks_29_ce1),
        .cnt_bucket_chunks_29_d1(cnt_bucket_chunks_29_d1),
        .cnt_bucket_chunks_29_q1(cnt_bucket_chunks_29_q1),
        .cnt_bucket_chunks_29_we1(cnt_bucket_chunks_29_we1),
        .cnt_bucket_chunks_30_address0(cnt_bucket_chunks_30_address0),
        .cnt_bucket_chunks_30_ce0(cnt_bucket_chunks_30_ce0),
        .cnt_bucket_chunks_30_d0(cnt_bucket_chunks_30_d0),
        .cnt_bucket_chunks_30_q0(cnt_bucket_chunks_30_q0),
        .cnt_bucket_chunks_30_we0(cnt_bucket_chunks_30_we0),
        .cnt_bucket_chunks_30_address1(cnt_bucket_chunks_30_address1),
        .cnt_bucket_chunks_30_ce1(cnt_bucket_chunks_30_ce1),
        .cnt_bucket_chunks_30_d1(cnt_bucket_chunks_30_d1),
        .cnt_bucket_chunks_30_q1(cnt_bucket_chunks_30_q1),
        .cnt_bucket_chunks_30_we1(cnt_bucket_chunks_30_we1),
        .cnt_bucket_chunks_31_address0(cnt_bucket_chunks_31_address0),
        .cnt_bucket_chunks_31_ce0(cnt_bucket_chunks_31_ce0),
        .cnt_bucket_chunks_31_d0(cnt_bucket_chunks_31_d0),
        .cnt_bucket_chunks_31_q0(cnt_bucket_chunks_31_q0),
        .cnt_bucket_chunks_31_we0(cnt_bucket_chunks_31_we0),
        .cnt_bucket_chunks_31_address1(cnt_bucket_chunks_31_address1),
        .cnt_bucket_chunks_31_ce1(cnt_bucket_chunks_31_ce1),
        .cnt_bucket_chunks_31_d1(cnt_bucket_chunks_31_d1),
        .cnt_bucket_chunks_31_q1(cnt_bucket_chunks_31_q1),
        .cnt_bucket_chunks_31_we1(cnt_bucket_chunks_31_we1),
        .cnt_bucket_chunks_32_address0(cnt_bucket_chunks_32_address0),
        .cnt_bucket_chunks_32_ce0(cnt_bucket_chunks_32_ce0),
        .cnt_bucket_chunks_32_d0(cnt_bucket_chunks_32_d0),
        .cnt_bucket_chunks_32_q0(cnt_bucket_chunks_32_q0),
        .cnt_bucket_chunks_32_we0(cnt_bucket_chunks_32_we0),
        .cnt_bucket_chunks_32_address1(cnt_bucket_chunks_32_address1),
        .cnt_bucket_chunks_32_ce1(cnt_bucket_chunks_32_ce1),
        .cnt_bucket_chunks_32_d1(cnt_bucket_chunks_32_d1),
        .cnt_bucket_chunks_32_q1(cnt_bucket_chunks_32_q1),
        .cnt_bucket_chunks_32_we1(cnt_bucket_chunks_32_we1),
        .cnt_bucket_chunks_33_address0(cnt_bucket_chunks_33_address0),
        .cnt_bucket_chunks_33_ce0(cnt_bucket_chunks_33_ce0),
        .cnt_bucket_chunks_33_d0(cnt_bucket_chunks_33_d0),
        .cnt_bucket_chunks_33_q0(cnt_bucket_chunks_33_q0),
        .cnt_bucket_chunks_33_we0(cnt_bucket_chunks_33_we0),
        .cnt_bucket_chunks_33_address1(cnt_bucket_chunks_33_address1),
        .cnt_bucket_chunks_33_ce1(cnt_bucket_chunks_33_ce1),
        .cnt_bucket_chunks_33_d1(cnt_bucket_chunks_33_d1),
        .cnt_bucket_chunks_33_q1(cnt_bucket_chunks_33_q1),
        .cnt_bucket_chunks_33_we1(cnt_bucket_chunks_33_we1),
        .cnt_bucket_chunks_34_address0(cnt_bucket_chunks_34_address0),
        .cnt_bucket_chunks_34_ce0(cnt_bucket_chunks_34_ce0),
        .cnt_bucket_chunks_34_d0(cnt_bucket_chunks_34_d0),
        .cnt_bucket_chunks_34_q0(cnt_bucket_chunks_34_q0),
        .cnt_bucket_chunks_34_we0(cnt_bucket_chunks_34_we0),
        .cnt_bucket_chunks_34_address1(cnt_bucket_chunks_34_address1),
        .cnt_bucket_chunks_34_ce1(cnt_bucket_chunks_34_ce1),
        .cnt_bucket_chunks_34_d1(cnt_bucket_chunks_34_d1),
        .cnt_bucket_chunks_34_q1(cnt_bucket_chunks_34_q1),
        .cnt_bucket_chunks_34_we1(cnt_bucket_chunks_34_we1),
        .cnt_bucket_chunks_35_address0(cnt_bucket_chunks_35_address0),
        .cnt_bucket_chunks_35_ce0(cnt_bucket_chunks_35_ce0),
        .cnt_bucket_chunks_35_d0(cnt_bucket_chunks_35_d0),
        .cnt_bucket_chunks_35_q0(cnt_bucket_chunks_35_q0),
        .cnt_bucket_chunks_35_we0(cnt_bucket_chunks_35_we0),
        .cnt_bucket_chunks_35_address1(cnt_bucket_chunks_35_address1),
        .cnt_bucket_chunks_35_ce1(cnt_bucket_chunks_35_ce1),
        .cnt_bucket_chunks_35_d1(cnt_bucket_chunks_35_d1),
        .cnt_bucket_chunks_35_q1(cnt_bucket_chunks_35_q1),
        .cnt_bucket_chunks_35_we1(cnt_bucket_chunks_35_we1),
        .cnt_bucket_chunks_36_address0(cnt_bucket_chunks_36_address0),
        .cnt_bucket_chunks_36_ce0(cnt_bucket_chunks_36_ce0),
        .cnt_bucket_chunks_36_d0(cnt_bucket_chunks_36_d0),
        .cnt_bucket_chunks_36_q0(cnt_bucket_chunks_36_q0),
        .cnt_bucket_chunks_36_we0(cnt_bucket_chunks_36_we0),
        .cnt_bucket_chunks_36_address1(cnt_bucket_chunks_36_address1),
        .cnt_bucket_chunks_36_ce1(cnt_bucket_chunks_36_ce1),
        .cnt_bucket_chunks_36_d1(cnt_bucket_chunks_36_d1),
        .cnt_bucket_chunks_36_q1(cnt_bucket_chunks_36_q1),
        .cnt_bucket_chunks_36_we1(cnt_bucket_chunks_36_we1),
        .cnt_bucket_chunks_37_address0(cnt_bucket_chunks_37_address0),
        .cnt_bucket_chunks_37_ce0(cnt_bucket_chunks_37_ce0),
        .cnt_bucket_chunks_37_d0(cnt_bucket_chunks_37_d0),
        .cnt_bucket_chunks_37_q0(cnt_bucket_chunks_37_q0),
        .cnt_bucket_chunks_37_we0(cnt_bucket_chunks_37_we0),
        .cnt_bucket_chunks_37_address1(cnt_bucket_chunks_37_address1),
        .cnt_bucket_chunks_37_ce1(cnt_bucket_chunks_37_ce1),
        .cnt_bucket_chunks_37_d1(cnt_bucket_chunks_37_d1),
        .cnt_bucket_chunks_37_q1(cnt_bucket_chunks_37_q1),
        .cnt_bucket_chunks_37_we1(cnt_bucket_chunks_37_we1),
        .cnt_bucket_chunks_38_address0(cnt_bucket_chunks_38_address0),
        .cnt_bucket_chunks_38_ce0(cnt_bucket_chunks_38_ce0),
        .cnt_bucket_chunks_38_d0(cnt_bucket_chunks_38_d0),
        .cnt_bucket_chunks_38_q0(cnt_bucket_chunks_38_q0),
        .cnt_bucket_chunks_38_we0(cnt_bucket_chunks_38_we0),
        .cnt_bucket_chunks_38_address1(cnt_bucket_chunks_38_address1),
        .cnt_bucket_chunks_38_ce1(cnt_bucket_chunks_38_ce1),
        .cnt_bucket_chunks_38_d1(cnt_bucket_chunks_38_d1),
        .cnt_bucket_chunks_38_q1(cnt_bucket_chunks_38_q1),
        .cnt_bucket_chunks_38_we1(cnt_bucket_chunks_38_we1),
        .cnt_bucket_chunks_39_address0(cnt_bucket_chunks_39_address0),
        .cnt_bucket_chunks_39_ce0(cnt_bucket_chunks_39_ce0),
        .cnt_bucket_chunks_39_d0(cnt_bucket_chunks_39_d0),
        .cnt_bucket_chunks_39_q0(cnt_bucket_chunks_39_q0),
        .cnt_bucket_chunks_39_we0(cnt_bucket_chunks_39_we0),
        .cnt_bucket_chunks_39_address1(cnt_bucket_chunks_39_address1),
        .cnt_bucket_chunks_39_ce1(cnt_bucket_chunks_39_ce1),
        .cnt_bucket_chunks_39_d1(cnt_bucket_chunks_39_d1),
        .cnt_bucket_chunks_39_q1(cnt_bucket_chunks_39_q1),
        .cnt_bucket_chunks_39_we1(cnt_bucket_chunks_39_we1),
        .cnt_bucket_chunks_40_address0(cnt_bucket_chunks_40_address0),
        .cnt_bucket_chunks_40_ce0(cnt_bucket_chunks_40_ce0),
        .cnt_bucket_chunks_40_d0(cnt_bucket_chunks_40_d0),
        .cnt_bucket_chunks_40_q0(cnt_bucket_chunks_40_q0),
        .cnt_bucket_chunks_40_we0(cnt_bucket_chunks_40_we0),
        .cnt_bucket_chunks_40_address1(cnt_bucket_chunks_40_address1),
        .cnt_bucket_chunks_40_ce1(cnt_bucket_chunks_40_ce1),
        .cnt_bucket_chunks_40_d1(cnt_bucket_chunks_40_d1),
        .cnt_bucket_chunks_40_q1(cnt_bucket_chunks_40_q1),
        .cnt_bucket_chunks_40_we1(cnt_bucket_chunks_40_we1),
        .cnt_bucket_chunks_41_address0(cnt_bucket_chunks_41_address0),
        .cnt_bucket_chunks_41_ce0(cnt_bucket_chunks_41_ce0),
        .cnt_bucket_chunks_41_d0(cnt_bucket_chunks_41_d0),
        .cnt_bucket_chunks_41_q0(cnt_bucket_chunks_41_q0),
        .cnt_bucket_chunks_41_we0(cnt_bucket_chunks_41_we0),
        .cnt_bucket_chunks_41_address1(cnt_bucket_chunks_41_address1),
        .cnt_bucket_chunks_41_ce1(cnt_bucket_chunks_41_ce1),
        .cnt_bucket_chunks_41_d1(cnt_bucket_chunks_41_d1),
        .cnt_bucket_chunks_41_q1(cnt_bucket_chunks_41_q1),
        .cnt_bucket_chunks_41_we1(cnt_bucket_chunks_41_we1),
        .cnt_bucket_chunks_42_address0(cnt_bucket_chunks_42_address0),
        .cnt_bucket_chunks_42_ce0(cnt_bucket_chunks_42_ce0),
        .cnt_bucket_chunks_42_d0(cnt_bucket_chunks_42_d0),
        .cnt_bucket_chunks_42_q0(cnt_bucket_chunks_42_q0),
        .cnt_bucket_chunks_42_we0(cnt_bucket_chunks_42_we0),
        .cnt_bucket_chunks_42_address1(cnt_bucket_chunks_42_address1),
        .cnt_bucket_chunks_42_ce1(cnt_bucket_chunks_42_ce1),
        .cnt_bucket_chunks_42_d1(cnt_bucket_chunks_42_d1),
        .cnt_bucket_chunks_42_q1(cnt_bucket_chunks_42_q1),
        .cnt_bucket_chunks_42_we1(cnt_bucket_chunks_42_we1),
        .num_padd_ops_dout(num_padd_ops_test_mem_data),
        .num_padd_ops_empty_n(num_padd_ops_stream_empty_n),
        .num_padd_ops_read(num_padd_ops_stream_read),
        .total_num_padd_ops(total_num_padd_ops)
        // .ap_return(msm_return)
    );

    test_case_memory  #( .EC_BASE_FIELD_WIDTH(EC_BASE_FIELD_WIDTH), .EC_SCALAR_FIELD_WIDTH(EC_SCALAR_FIELD_WIDTH), .ADDR_WIDTH(ADDR_WIDTH), .MEM_SIZE(MEM_SIZE)) test_case_mem_0 (
        ap_clk, ap_rst, debug, 
        P_arr_x_address0, P_arr_x_ce0, P_arr_x_d0, P_arr_x_q0, P_arr_x_we0,
        P_arr_x_address1, P_arr_x_ce1, P_arr_x_d1, P_arr_x_q1, P_arr_x_we1,
        P_arr_y_address0, P_arr_y_ce0, P_arr_y_d0, P_arr_y_q0, P_arr_y_we0,
        P_arr_y_address1, P_arr_y_ce1, P_arr_y_d1, P_arr_y_q1, P_arr_y_we1,
        P_arr_z_address0, P_arr_z_ce0, P_arr_z_d0, P_arr_z_q0, P_arr_z_we0,
        P_arr_z_address1, P_arr_z_ce1, P_arr_z_d1, P_arr_z_q1, P_arr_z_we1,
        K_arr_address0, K_arr_ce0, K_arr_d0, K_arr_q0, K_arr_we0,
        K_arr_address1, K_arr_ce1, K_arr_d1, K_arr_q1, K_arr_we1,
        total_num_padd_ops, read_count, count_test_mem_data, read_num_padd_ops,
        num_padd_ops_test_mem_data,
        B_i_address0, B_i_ce0, B_i_d0, B_i_q0, B_i_we0, B_i_address1, B_i_ce1, B_i_d1, B_i_q1, B_i_we1
    );

endmodule
